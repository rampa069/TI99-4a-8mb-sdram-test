
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c4",x"ee",x"c2"),
    14 => (x"48",x"e8",x"da",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e9",x"e2"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"e8",x"da"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"da",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"e8"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"ec",x"da",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"f0",x"da",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"f0",x"da",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"f0",x"da"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"f7",x"da"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"f8",x"da"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"f9",x"da",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"da",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"f9"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"fa",x"da",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"f5",x"da"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"f6",x"da",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"da",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"f7"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"f8",x"da",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e3",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"d6"),
   330 => (x"1e",x"ce",x"db",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"e2",x"f2",x"c0",x"7e"),
   337 => (x"dc",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"c4"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"de",x"f2"),
   343 => (x"4a",x"e0",x"dc",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e2",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"d4"),
   350 => (x"bf",x"9f",x"cc",x"e3"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"d4",x"e2",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"db",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"ce"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"de",x"f2"),
   365 => (x"4a",x"e0",x"dc",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"d6",x"e3"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"e2",x"f2"),
   372 => (x"4a",x"c4",x"dc",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"cc",x"e3",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e3",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"cd"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"ce",x"db",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"d9",x"db",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"da",x"db"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"db",x"db",x"c2"),
   400 => (x"e3",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"d2"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"d6",x"e3"),
   404 => (x"bf",x"97",x"dc",x"db"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"dd",x"db"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e7",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"e3"),
   410 => (x"97",x"de",x"db",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"d6",x"e3",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"de",x"f2",x"c0",x"87"),
   415 => (x"dc",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"e0"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"ce",x"e3"),
   422 => (x"5c",x"f7",x"e7",x"c2"),
   423 => (x"97",x"f3",x"db",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"f2",x"db",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"f4",x"db",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"f5",x"db"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"e3",x"e7",x"c2",x"91"),
   434 => (x"e7",x"c2",x"81",x"bf"),
   435 => (x"db",x"c2",x"59",x"eb"),
   436 => (x"4a",x"bf",x"97",x"fb"),
   437 => (x"db",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"fa"),
   439 => (x"db",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"fc"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"fd",x"db",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e7",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"ef"),
   447 => (x"e7",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"ef"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"e0",x"db",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"df",x"db",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"f7",x"e7"),
   457 => (x"bf",x"97",x"e5",x"db"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"e4",x"db"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"f3",x"e7",x"c2"),
   463 => (x"48",x"eb",x"e7",x"c2"),
   464 => (x"e7",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"e7"),
   466 => (x"f7",x"e7",x"c2",x"78"),
   467 => (x"eb",x"e7",x"c2",x"48"),
   468 => (x"e7",x"c2",x"78",x"bf"),
   469 => (x"e7",x"c2",x"48",x"fb"),
   470 => (x"c2",x"78",x"bf",x"ef"),
   471 => (x"02",x"bf",x"d6",x"e3"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"f3",x"e7",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"da",x"e3",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"d6",x"e3"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e7",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"e3"),
   492 => (x"ab",x"bf",x"da",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"de",x"f2"),
   495 => (x"73",x"1e",x"ce",x"db"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"d6",x"e3",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"ce",x"db"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"ce",x"db",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c1",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"ea",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d6",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"de",x"e3",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d4",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"cf",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"d6",x"e3"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"49",x"6e",x"7e",x"c0"),
   556 => (x"bf",x"66",x"c4",x"48"),
   557 => (x"08",x"66",x"c4",x"80"),
   558 => (x"cc",x"7c",x"c0",x"78"),
   559 => (x"66",x"c4",x"49",x"a4"),
   560 => (x"a4",x"d0",x"79",x"bf"),
   561 => (x"c1",x"79",x"c0",x"49"),
   562 => (x"c0",x"87",x"c2",x"48"),
   563 => (x"fa",x"8e",x"f8",x"48"),
   564 => (x"5e",x"0e",x"87",x"ed"),
   565 => (x"0e",x"5d",x"5c",x"5b"),
   566 => (x"02",x"9c",x"4c",x"71"),
   567 => (x"c8",x"87",x"cb",x"c1"),
   568 => (x"02",x"69",x"49",x"a4"),
   569 => (x"d0",x"87",x"c3",x"c1"),
   570 => (x"49",x"6c",x"4a",x"66"),
   571 => (x"72",x"48",x"a6",x"d0"),
   572 => (x"b9",x"4d",x"78",x"a1"),
   573 => (x"bf",x"d2",x"e3",x"c2"),
   574 => (x"72",x"ba",x"ff",x"4a"),
   575 => (x"02",x"99",x"71",x"99"),
   576 => (x"c4",x"87",x"e4",x"c0"),
   577 => (x"49",x"6b",x"4b",x"a4"),
   578 => (x"70",x"87",x"fc",x"f9"),
   579 => (x"ce",x"e3",x"c2",x"7b"),
   580 => (x"81",x"6c",x"49",x"bf"),
   581 => (x"b9",x"75",x"7c",x"71"),
   582 => (x"bf",x"d2",x"e3",x"c2"),
   583 => (x"72",x"ba",x"ff",x"4a"),
   584 => (x"05",x"99",x"71",x"99"),
   585 => (x"d0",x"87",x"dc",x"ff"),
   586 => (x"d2",x"f9",x"7c",x"66"),
   587 => (x"1e",x"73",x"1e",x"87"),
   588 => (x"02",x"9b",x"4b",x"71"),
   589 => (x"a3",x"c8",x"87",x"c7"),
   590 => (x"c5",x"05",x"69",x"49"),
   591 => (x"c0",x"48",x"c0",x"87"),
   592 => (x"e7",x"c2",x"87",x"f6"),
   593 => (x"c4",x"49",x"bf",x"e7"),
   594 => (x"4a",x"6a",x"4a",x"a3"),
   595 => (x"e3",x"c2",x"8a",x"c2"),
   596 => (x"72",x"92",x"bf",x"ce"),
   597 => (x"e3",x"c2",x"49",x"a1"),
   598 => (x"6b",x"4a",x"bf",x"d2"),
   599 => (x"49",x"a1",x"72",x"9a"),
   600 => (x"59",x"de",x"f2",x"c0"),
   601 => (x"71",x"1e",x"66",x"c8"),
   602 => (x"c4",x"87",x"e4",x"ea"),
   603 => (x"05",x"98",x"70",x"86"),
   604 => (x"48",x"c0",x"87",x"c4"),
   605 => (x"48",x"c1",x"87",x"c2"),
   606 => (x"1e",x"87",x"c8",x"f8"),
   607 => (x"4b",x"71",x"1e",x"73"),
   608 => (x"87",x"c7",x"02",x"9b"),
   609 => (x"69",x"49",x"a3",x"c8"),
   610 => (x"c0",x"87",x"c5",x"05"),
   611 => (x"87",x"f6",x"c0",x"48"),
   612 => (x"bf",x"e7",x"e7",x"c2"),
   613 => (x"4a",x"a3",x"c4",x"49"),
   614 => (x"8a",x"c2",x"4a",x"6a"),
   615 => (x"bf",x"ce",x"e3",x"c2"),
   616 => (x"49",x"a1",x"72",x"92"),
   617 => (x"bf",x"d2",x"e3",x"c2"),
   618 => (x"72",x"9a",x"6b",x"4a"),
   619 => (x"f2",x"c0",x"49",x"a1"),
   620 => (x"66",x"c8",x"59",x"de"),
   621 => (x"cf",x"e6",x"71",x"1e"),
   622 => (x"70",x"86",x"c4",x"87"),
   623 => (x"87",x"c4",x"05",x"98"),
   624 => (x"87",x"c2",x"48",x"c0"),
   625 => (x"fa",x"f6",x"48",x"c1"),
   626 => (x"5b",x"5e",x"0e",x"87"),
   627 => (x"1e",x"0e",x"5d",x"5c"),
   628 => (x"66",x"d4",x"4b",x"71"),
   629 => (x"02",x"9b",x"73",x"4d"),
   630 => (x"c8",x"87",x"cc",x"c1"),
   631 => (x"02",x"69",x"49",x"a3"),
   632 => (x"d0",x"87",x"c4",x"c1"),
   633 => (x"e3",x"c2",x"4c",x"a3"),
   634 => (x"ff",x"49",x"bf",x"d2"),
   635 => (x"99",x"4a",x"6c",x"b9"),
   636 => (x"a9",x"66",x"d4",x"7e"),
   637 => (x"c0",x"87",x"cd",x"06"),
   638 => (x"a3",x"cc",x"7c",x"7b"),
   639 => (x"49",x"a3",x"c4",x"4a"),
   640 => (x"87",x"ca",x"79",x"6a"),
   641 => (x"c0",x"f8",x"49",x"72"),
   642 => (x"4d",x"66",x"d4",x"99"),
   643 => (x"49",x"75",x"8d",x"71"),
   644 => (x"1e",x"71",x"29",x"c9"),
   645 => (x"f9",x"fa",x"49",x"73"),
   646 => (x"ce",x"db",x"c2",x"87"),
   647 => (x"fc",x"49",x"73",x"1e"),
   648 => (x"86",x"c8",x"87",x"cb"),
   649 => (x"26",x"7c",x"66",x"d4"),
   650 => (x"1e",x"87",x"d4",x"f5"),
   651 => (x"4b",x"71",x"1e",x"73"),
   652 => (x"e4",x"c0",x"02",x"9b"),
   653 => (x"fb",x"e7",x"c2",x"87"),
   654 => (x"c2",x"4a",x"73",x"5b"),
   655 => (x"ce",x"e3",x"c2",x"8a"),
   656 => (x"c2",x"92",x"49",x"bf"),
   657 => (x"48",x"bf",x"e7",x"e7"),
   658 => (x"e7",x"c2",x"80",x"72"),
   659 => (x"48",x"71",x"58",x"ff"),
   660 => (x"e3",x"c2",x"30",x"c4"),
   661 => (x"ed",x"c0",x"58",x"de"),
   662 => (x"f7",x"e7",x"c2",x"87"),
   663 => (x"eb",x"e7",x"c2",x"48"),
   664 => (x"e7",x"c2",x"78",x"bf"),
   665 => (x"e7",x"c2",x"48",x"fb"),
   666 => (x"c2",x"78",x"bf",x"ef"),
   667 => (x"02",x"bf",x"d6",x"e3"),
   668 => (x"e3",x"c2",x"87",x"c9"),
   669 => (x"c4",x"49",x"bf",x"ce"),
   670 => (x"c2",x"87",x"c7",x"31"),
   671 => (x"49",x"bf",x"f3",x"e7"),
   672 => (x"e3",x"c2",x"31",x"c4"),
   673 => (x"fa",x"f3",x"59",x"de"),
   674 => (x"5b",x"5e",x"0e",x"87"),
   675 => (x"4a",x"71",x"0e",x"5c"),
   676 => (x"9a",x"72",x"4b",x"c0"),
   677 => (x"87",x"e1",x"c0",x"02"),
   678 => (x"9f",x"49",x"a2",x"da"),
   679 => (x"e3",x"c2",x"4b",x"69"),
   680 => (x"cf",x"02",x"bf",x"d6"),
   681 => (x"49",x"a2",x"d4",x"87"),
   682 => (x"4c",x"49",x"69",x"9f"),
   683 => (x"9c",x"ff",x"ff",x"c0"),
   684 => (x"87",x"c2",x"34",x"d0"),
   685 => (x"49",x"74",x"4c",x"c0"),
   686 => (x"fd",x"49",x"73",x"b3"),
   687 => (x"c0",x"f3",x"87",x"ed"),
   688 => (x"5b",x"5e",x"0e",x"87"),
   689 => (x"f4",x"0e",x"5d",x"5c"),
   690 => (x"c0",x"4a",x"71",x"86"),
   691 => (x"02",x"9a",x"72",x"7e"),
   692 => (x"db",x"c2",x"87",x"d8"),
   693 => (x"78",x"c0",x"48",x"ca"),
   694 => (x"48",x"c2",x"db",x"c2"),
   695 => (x"bf",x"fb",x"e7",x"c2"),
   696 => (x"c6",x"db",x"c2",x"78"),
   697 => (x"f7",x"e7",x"c2",x"48"),
   698 => (x"e3",x"c2",x"78",x"bf"),
   699 => (x"50",x"c0",x"48",x"eb"),
   700 => (x"bf",x"da",x"e3",x"c2"),
   701 => (x"ca",x"db",x"c2",x"49"),
   702 => (x"aa",x"71",x"4a",x"bf"),
   703 => (x"87",x"c9",x"c4",x"03"),
   704 => (x"99",x"cf",x"49",x"72"),
   705 => (x"87",x"e9",x"c0",x"05"),
   706 => (x"48",x"da",x"f2",x"c0"),
   707 => (x"bf",x"c2",x"db",x"c2"),
   708 => (x"ce",x"db",x"c2",x"78"),
   709 => (x"c2",x"db",x"c2",x"1e"),
   710 => (x"db",x"c2",x"49",x"bf"),
   711 => (x"a1",x"c1",x"48",x"c2"),
   712 => (x"ea",x"e3",x"71",x"78"),
   713 => (x"c0",x"86",x"c4",x"87"),
   714 => (x"c2",x"48",x"d6",x"f2"),
   715 => (x"cc",x"78",x"ce",x"db"),
   716 => (x"d6",x"f2",x"c0",x"87"),
   717 => (x"e0",x"c0",x"48",x"bf"),
   718 => (x"da",x"f2",x"c0",x"80"),
   719 => (x"ca",x"db",x"c2",x"58"),
   720 => (x"80",x"c1",x"48",x"bf"),
   721 => (x"58",x"ce",x"db",x"c2"),
   722 => (x"00",x"0c",x"96",x"27"),
   723 => (x"bf",x"97",x"bf",x"00"),
   724 => (x"c2",x"02",x"9d",x"4d"),
   725 => (x"e5",x"c3",x"87",x"e3"),
   726 => (x"dc",x"c2",x"02",x"ad"),
   727 => (x"d6",x"f2",x"c0",x"87"),
   728 => (x"a3",x"cb",x"4b",x"bf"),
   729 => (x"cf",x"4c",x"11",x"49"),
   730 => (x"d2",x"c1",x"05",x"ac"),
   731 => (x"df",x"49",x"75",x"87"),
   732 => (x"cd",x"89",x"c1",x"99"),
   733 => (x"de",x"e3",x"c2",x"91"),
   734 => (x"4a",x"a3",x"c1",x"81"),
   735 => (x"a3",x"c3",x"51",x"12"),
   736 => (x"c5",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"c7"),
   739 => (x"4a",x"a3",x"c9",x"51"),
   740 => (x"a3",x"ce",x"51",x"12"),
   741 => (x"d0",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"12",x"4a",x"a3",x"d2"),
   744 => (x"4a",x"a3",x"d4",x"51"),
   745 => (x"a3",x"d6",x"51",x"12"),
   746 => (x"d8",x"51",x"12",x"4a"),
   747 => (x"51",x"12",x"4a",x"a3"),
   748 => (x"12",x"4a",x"a3",x"dc"),
   749 => (x"4a",x"a3",x"de",x"51"),
   750 => (x"7e",x"c1",x"51",x"12"),
   751 => (x"74",x"87",x"fa",x"c0"),
   752 => (x"05",x"99",x"c8",x"49"),
   753 => (x"74",x"87",x"eb",x"c0"),
   754 => (x"05",x"99",x"d0",x"49"),
   755 => (x"66",x"dc",x"87",x"d1"),
   756 => (x"87",x"cb",x"c0",x"02"),
   757 => (x"66",x"dc",x"49",x"73"),
   758 => (x"02",x"98",x"70",x"0f"),
   759 => (x"6e",x"87",x"d3",x"c0"),
   760 => (x"87",x"c6",x"c0",x"05"),
   761 => (x"48",x"de",x"e3",x"c2"),
   762 => (x"f2",x"c0",x"50",x"c0"),
   763 => (x"c2",x"48",x"bf",x"d6"),
   764 => (x"e3",x"c2",x"87",x"df"),
   765 => (x"50",x"c0",x"48",x"eb"),
   766 => (x"da",x"e3",x"c2",x"7e"),
   767 => (x"db",x"c2",x"49",x"bf"),
   768 => (x"71",x"4a",x"bf",x"ca"),
   769 => (x"f7",x"fb",x"04",x"aa"),
   770 => (x"fb",x"e7",x"c2",x"87"),
   771 => (x"c8",x"c0",x"05",x"bf"),
   772 => (x"d6",x"e3",x"c2",x"87"),
   773 => (x"f6",x"c1",x"02",x"bf"),
   774 => (x"c6",x"db",x"c2",x"87"),
   775 => (x"e6",x"ed",x"49",x"bf"),
   776 => (x"ca",x"db",x"c2",x"87"),
   777 => (x"48",x"a6",x"c4",x"58"),
   778 => (x"bf",x"c6",x"db",x"c2"),
   779 => (x"d6",x"e3",x"c2",x"78"),
   780 => (x"d8",x"c0",x"02",x"bf"),
   781 => (x"49",x"66",x"c4",x"87"),
   782 => (x"ff",x"ff",x"ff",x"cf"),
   783 => (x"02",x"a9",x"99",x"f8"),
   784 => (x"c0",x"87",x"c5",x"c0"),
   785 => (x"87",x"e1",x"c0",x"4c"),
   786 => (x"dc",x"c0",x"4c",x"c1"),
   787 => (x"49",x"66",x"c4",x"87"),
   788 => (x"99",x"f8",x"ff",x"cf"),
   789 => (x"c8",x"c0",x"02",x"a9"),
   790 => (x"48",x"a6",x"c8",x"87"),
   791 => (x"c5",x"c0",x"78",x"c0"),
   792 => (x"48",x"a6",x"c8",x"87"),
   793 => (x"66",x"c8",x"78",x"c1"),
   794 => (x"05",x"9c",x"74",x"4c"),
   795 => (x"c4",x"87",x"e0",x"c0"),
   796 => (x"89",x"c2",x"49",x"66"),
   797 => (x"bf",x"ce",x"e3",x"c2"),
   798 => (x"e7",x"c2",x"91",x"4a"),
   799 => (x"c2",x"4a",x"bf",x"e7"),
   800 => (x"72",x"48",x"c2",x"db"),
   801 => (x"db",x"c2",x"78",x"a1"),
   802 => (x"78",x"c0",x"48",x"ca"),
   803 => (x"c0",x"87",x"e1",x"f9"),
   804 => (x"eb",x"8e",x"f4",x"48"),
   805 => (x"00",x"00",x"87",x"e9"),
   806 => (x"ff",x"ff",x"00",x"00"),
   807 => (x"0c",x"a6",x"ff",x"ff"),
   808 => (x"0c",x"af",x"00",x"00"),
   809 => (x"41",x"46",x"00",x"00"),
   810 => (x"20",x"32",x"33",x"54"),
   811 => (x"46",x"00",x"20",x"20"),
   812 => (x"36",x"31",x"54",x"41"),
   813 => (x"00",x"20",x"20",x"20"),
   814 => (x"48",x"d4",x"ff",x"1e"),
   815 => (x"68",x"78",x"ff",x"c3"),
   816 => (x"1e",x"4f",x"26",x"48"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"d0",x"ff",x"78",x"ff"),
   819 => (x"78",x"e1",x"c0",x"48"),
   820 => (x"d4",x"48",x"d4",x"ff"),
   821 => (x"ff",x"e7",x"c2",x"78"),
   822 => (x"bf",x"d4",x"ff",x"48"),
   823 => (x"1e",x"4f",x"26",x"50"),
   824 => (x"c0",x"48",x"d0",x"ff"),
   825 => (x"4f",x"26",x"78",x"e0"),
   826 => (x"87",x"cc",x"ff",x"1e"),
   827 => (x"02",x"99",x"49",x"70"),
   828 => (x"fb",x"c0",x"87",x"c6"),
   829 => (x"87",x"f1",x"05",x"a9"),
   830 => (x"4f",x"26",x"48",x"71"),
   831 => (x"5c",x"5b",x"5e",x"0e"),
   832 => (x"c0",x"4b",x"71",x"0e"),
   833 => (x"87",x"f0",x"fe",x"4c"),
   834 => (x"02",x"99",x"49",x"70"),
   835 => (x"c0",x"87",x"f9",x"c0"),
   836 => (x"c0",x"02",x"a9",x"ec"),
   837 => (x"fb",x"c0",x"87",x"f2"),
   838 => (x"eb",x"c0",x"02",x"a9"),
   839 => (x"b7",x"66",x"cc",x"87"),
   840 => (x"87",x"c7",x"03",x"ac"),
   841 => (x"c2",x"02",x"66",x"d0"),
   842 => (x"71",x"53",x"71",x"87"),
   843 => (x"87",x"c2",x"02",x"99"),
   844 => (x"c3",x"fe",x"84",x"c1"),
   845 => (x"99",x"49",x"70",x"87"),
   846 => (x"c0",x"87",x"cd",x"02"),
   847 => (x"c7",x"02",x"a9",x"ec"),
   848 => (x"a9",x"fb",x"c0",x"87"),
   849 => (x"87",x"d5",x"ff",x"05"),
   850 => (x"c3",x"02",x"66",x"d0"),
   851 => (x"7b",x"97",x"c0",x"87"),
   852 => (x"05",x"a9",x"ec",x"c0"),
   853 => (x"4a",x"74",x"87",x"c4"),
   854 => (x"4a",x"74",x"87",x"c5"),
   855 => (x"72",x"8a",x"0a",x"c0"),
   856 => (x"26",x"87",x"c2",x"48"),
   857 => (x"26",x"4c",x"26",x"4d"),
   858 => (x"1e",x"4f",x"26",x"4b"),
   859 => (x"70",x"87",x"c9",x"fd"),
   860 => (x"aa",x"f0",x"c0",x"4a"),
   861 => (x"c0",x"87",x"c9",x"04"),
   862 => (x"c3",x"01",x"aa",x"f9"),
   863 => (x"8a",x"f0",x"c0",x"87"),
   864 => (x"04",x"aa",x"c1",x"c1"),
   865 => (x"da",x"c1",x"87",x"c9"),
   866 => (x"87",x"c3",x"01",x"aa"),
   867 => (x"72",x"8a",x"f7",x"c0"),
   868 => (x"0e",x"4f",x"26",x"48"),
   869 => (x"5d",x"5c",x"5b",x"5e"),
   870 => (x"71",x"86",x"f8",x"0e"),
   871 => (x"fc",x"7e",x"c0",x"4c"),
   872 => (x"4b",x"c0",x"87",x"e1"),
   873 => (x"97",x"c0",x"f9",x"c0"),
   874 => (x"a9",x"c0",x"49",x"bf"),
   875 => (x"fc",x"87",x"cf",x"04"),
   876 => (x"83",x"c1",x"87",x"f6"),
   877 => (x"97",x"c0",x"f9",x"c0"),
   878 => (x"06",x"ab",x"49",x"bf"),
   879 => (x"f9",x"c0",x"87",x"f1"),
   880 => (x"02",x"bf",x"97",x"c0"),
   881 => (x"ef",x"fb",x"87",x"cf"),
   882 => (x"99",x"49",x"70",x"87"),
   883 => (x"c0",x"87",x"c6",x"02"),
   884 => (x"f1",x"05",x"a9",x"ec"),
   885 => (x"fb",x"4b",x"c0",x"87"),
   886 => (x"4d",x"70",x"87",x"de"),
   887 => (x"c8",x"87",x"d9",x"fb"),
   888 => (x"d3",x"fb",x"58",x"a6"),
   889 => (x"c1",x"4a",x"70",x"87"),
   890 => (x"49",x"a4",x"c8",x"83"),
   891 => (x"ad",x"49",x"69",x"97"),
   892 => (x"c0",x"87",x"c7",x"02"),
   893 => (x"c0",x"05",x"ad",x"ff"),
   894 => (x"a4",x"c9",x"87",x"e7"),
   895 => (x"49",x"69",x"97",x"49"),
   896 => (x"02",x"a9",x"66",x"c4"),
   897 => (x"c0",x"48",x"87",x"c7"),
   898 => (x"d4",x"05",x"a8",x"ff"),
   899 => (x"49",x"a4",x"ca",x"87"),
   900 => (x"aa",x"49",x"69",x"97"),
   901 => (x"c0",x"87",x"c6",x"02"),
   902 => (x"c4",x"05",x"aa",x"ff"),
   903 => (x"d0",x"7e",x"c1",x"87"),
   904 => (x"ad",x"ec",x"c0",x"87"),
   905 => (x"c0",x"87",x"c6",x"02"),
   906 => (x"c4",x"05",x"ad",x"fb"),
   907 => (x"c1",x"4b",x"c0",x"87"),
   908 => (x"fe",x"02",x"6e",x"7e"),
   909 => (x"e6",x"fa",x"87",x"e1"),
   910 => (x"f8",x"48",x"73",x"87"),
   911 => (x"87",x"e3",x"fc",x"8e"),
   912 => (x"5b",x"5e",x"0e",x"00"),
   913 => (x"f4",x"0e",x"5d",x"5c"),
   914 => (x"ff",x"7e",x"71",x"86"),
   915 => (x"1e",x"6e",x"4b",x"d4"),
   916 => (x"49",x"c4",x"e8",x"c2"),
   917 => (x"c4",x"87",x"e2",x"e6"),
   918 => (x"02",x"98",x"70",x"86"),
   919 => (x"c4",x"87",x"f5",x"c4"),
   920 => (x"e4",x"c1",x"48",x"a6"),
   921 => (x"6e",x"78",x"bf",x"cc"),
   922 => (x"87",x"e7",x"fc",x"49"),
   923 => (x"70",x"58",x"a6",x"cc"),
   924 => (x"87",x"c5",x"05",x"98"),
   925 => (x"c1",x"48",x"a6",x"c8"),
   926 => (x"48",x"d0",x"ff",x"78"),
   927 => (x"d5",x"c1",x"78",x"c5"),
   928 => (x"49",x"66",x"c8",x"7b"),
   929 => (x"31",x"c6",x"89",x"c1"),
   930 => (x"97",x"ca",x"e4",x"c1"),
   931 => (x"71",x"48",x"4a",x"bf"),
   932 => (x"ff",x"7b",x"70",x"b0"),
   933 => (x"78",x"c4",x"48",x"d0"),
   934 => (x"d6",x"c1",x"78",x"c5"),
   935 => (x"6e",x"4d",x"c0",x"7b"),
   936 => (x"11",x"81",x"75",x"49"),
   937 => (x"cb",x"85",x"c1",x"7b"),
   938 => (x"f2",x"04",x"ad",x"b7"),
   939 => (x"c3",x"4d",x"cc",x"87"),
   940 => (x"85",x"c1",x"7b",x"ff"),
   941 => (x"ad",x"b7",x"e0",x"c0"),
   942 => (x"ff",x"87",x"f4",x"04"),
   943 => (x"78",x"c4",x"48",x"d0"),
   944 => (x"c5",x"7b",x"ff",x"c3"),
   945 => (x"7b",x"d3",x"c1",x"78"),
   946 => (x"78",x"c4",x"7b",x"c1"),
   947 => (x"b7",x"c0",x"48",x"66"),
   948 => (x"ee",x"c2",x"06",x"a8"),
   949 => (x"cc",x"e8",x"c2",x"87"),
   950 => (x"66",x"c4",x"4c",x"bf"),
   951 => (x"c8",x"88",x"74",x"48"),
   952 => (x"9c",x"74",x"58",x"a6"),
   953 => (x"87",x"f7",x"c1",x"02"),
   954 => (x"7e",x"ce",x"db",x"c2"),
   955 => (x"8c",x"4d",x"c0",x"c8"),
   956 => (x"03",x"ac",x"b7",x"c0"),
   957 => (x"c0",x"c8",x"87",x"c6"),
   958 => (x"4c",x"c0",x"4d",x"a4"),
   959 => (x"97",x"ff",x"e7",x"c2"),
   960 => (x"99",x"d0",x"49",x"bf"),
   961 => (x"c0",x"87",x"d0",x"02"),
   962 => (x"c4",x"e8",x"c2",x"1e"),
   963 => (x"87",x"dd",x"e8",x"49"),
   964 => (x"4a",x"70",x"86",x"c4"),
   965 => (x"c2",x"87",x"ed",x"c0"),
   966 => (x"c2",x"1e",x"ce",x"db"),
   967 => (x"e8",x"49",x"c4",x"e8"),
   968 => (x"86",x"c4",x"87",x"cb"),
   969 => (x"d0",x"ff",x"4a",x"70"),
   970 => (x"78",x"c5",x"c8",x"48"),
   971 => (x"6e",x"7b",x"d4",x"c1"),
   972 => (x"6e",x"7b",x"bf",x"97"),
   973 => (x"70",x"80",x"c1",x"48"),
   974 => (x"05",x"8d",x"c1",x"7e"),
   975 => (x"ff",x"87",x"f0",x"ff"),
   976 => (x"78",x"c4",x"48",x"d0"),
   977 => (x"c5",x"05",x"9a",x"72"),
   978 => (x"c1",x"48",x"c0",x"87"),
   979 => (x"1e",x"c1",x"87",x"c8"),
   980 => (x"49",x"c4",x"e8",x"c2"),
   981 => (x"c4",x"87",x"fb",x"e5"),
   982 => (x"05",x"9c",x"74",x"86"),
   983 => (x"c4",x"87",x"c9",x"fe"),
   984 => (x"b7",x"c0",x"48",x"66"),
   985 => (x"87",x"d1",x"06",x"a8"),
   986 => (x"48",x"c4",x"e8",x"c2"),
   987 => (x"80",x"d0",x"78",x"c0"),
   988 => (x"80",x"f4",x"78",x"c0"),
   989 => (x"bf",x"d0",x"e8",x"c2"),
   990 => (x"48",x"66",x"c4",x"78"),
   991 => (x"01",x"a8",x"b7",x"c0"),
   992 => (x"ff",x"87",x"d2",x"fd"),
   993 => (x"78",x"c5",x"48",x"d0"),
   994 => (x"c0",x"7b",x"d3",x"c1"),
   995 => (x"c1",x"78",x"c4",x"7b"),
   996 => (x"87",x"c2",x"c0",x"48"),
   997 => (x"8e",x"f4",x"48",x"c0"),
   998 => (x"4c",x"26",x"4d",x"26"),
   999 => (x"4f",x"26",x"4b",x"26"),
  1000 => (x"5c",x"5b",x"5e",x"0e"),
  1001 => (x"71",x"1e",x"0e",x"5d"),
  1002 => (x"4d",x"4c",x"c0",x"4b"),
  1003 => (x"e8",x"c0",x"04",x"ab"),
  1004 => (x"d3",x"f6",x"c0",x"87"),
  1005 => (x"02",x"9d",x"75",x"1e"),
  1006 => (x"4a",x"c0",x"87",x"c4"),
  1007 => (x"4a",x"c1",x"87",x"c2"),
  1008 => (x"fc",x"eb",x"49",x"72"),
  1009 => (x"70",x"86",x"c4",x"87"),
  1010 => (x"6e",x"84",x"c1",x"7e"),
  1011 => (x"73",x"87",x"c2",x"05"),
  1012 => (x"73",x"85",x"c1",x"4c"),
  1013 => (x"d8",x"ff",x"06",x"ac"),
  1014 => (x"26",x"48",x"6e",x"87"),
  1015 => (x"0e",x"87",x"f9",x"fe"),
  1016 => (x"0e",x"5c",x"5b",x"5e"),
  1017 => (x"66",x"cc",x"4b",x"71"),
  1018 => (x"4c",x"87",x"d8",x"02"),
  1019 => (x"02",x"8c",x"f0",x"c0"),
  1020 => (x"4a",x"74",x"87",x"d8"),
  1021 => (x"d1",x"02",x"8a",x"c1"),
  1022 => (x"cd",x"02",x"8a",x"87"),
  1023 => (x"c9",x"02",x"8a",x"87"),
  1024 => (x"73",x"87",x"d9",x"87"),
  1025 => (x"87",x"f9",x"f8",x"49"),
  1026 => (x"1e",x"74",x"87",x"d2"),
  1027 => (x"d8",x"c1",x"49",x"c0"),
  1028 => (x"1e",x"74",x"87",x"d7"),
  1029 => (x"d8",x"c1",x"49",x"73"),
  1030 => (x"86",x"c8",x"87",x"cf"),
  1031 => (x"0e",x"87",x"fb",x"fd"),
  1032 => (x"5d",x"5c",x"5b",x"5e"),
  1033 => (x"4c",x"71",x"1e",x"0e"),
  1034 => (x"c2",x"91",x"de",x"49"),
  1035 => (x"71",x"4d",x"ec",x"e8"),
  1036 => (x"02",x"6d",x"97",x"85"),
  1037 => (x"c2",x"87",x"dc",x"c1"),
  1038 => (x"49",x"bf",x"d8",x"e8"),
  1039 => (x"fd",x"71",x"81",x"74"),
  1040 => (x"7e",x"70",x"87",x"de"),
  1041 => (x"c0",x"02",x"98",x"48"),
  1042 => (x"e8",x"c2",x"87",x"f2"),
  1043 => (x"4a",x"70",x"4b",x"e0"),
  1044 => (x"c1",x"ff",x"49",x"cb"),
  1045 => (x"4b",x"74",x"87",x"d1"),
  1046 => (x"e4",x"c1",x"93",x"cb"),
  1047 => (x"83",x"c4",x"83",x"de"),
  1048 => (x"7b",x"d7",x"c2",x"c1"),
  1049 => (x"c1",x"c1",x"49",x"74"),
  1050 => (x"7b",x"75",x"87",x"ed"),
  1051 => (x"97",x"cb",x"e4",x"c1"),
  1052 => (x"c2",x"1e",x"49",x"bf"),
  1053 => (x"fd",x"49",x"e0",x"e8"),
  1054 => (x"86",x"c4",x"87",x"e5"),
  1055 => (x"c1",x"c1",x"49",x"74"),
  1056 => (x"49",x"c0",x"87",x"d5"),
  1057 => (x"87",x"f4",x"c2",x"c1"),
  1058 => (x"48",x"c0",x"e8",x"c2"),
  1059 => (x"49",x"c1",x"78",x"c0"),
  1060 => (x"26",x"87",x"fb",x"dd"),
  1061 => (x"4c",x"87",x"c1",x"fc"),
  1062 => (x"69",x"64",x"61",x"6f"),
  1063 => (x"2e",x"2e",x"67",x"6e"),
  1064 => (x"73",x"1e",x"00",x"2e"),
  1065 => (x"49",x"4a",x"71",x"1e"),
  1066 => (x"bf",x"d8",x"e8",x"c2"),
  1067 => (x"ef",x"fb",x"71",x"81"),
  1068 => (x"9b",x"4b",x"70",x"87"),
  1069 => (x"49",x"87",x"c4",x"02"),
  1070 => (x"c2",x"87",x"ce",x"e7"),
  1071 => (x"c0",x"48",x"d8",x"e8"),
  1072 => (x"dd",x"49",x"c1",x"78"),
  1073 => (x"d3",x"fb",x"87",x"c8"),
  1074 => (x"49",x"c0",x"1e",x"87"),
  1075 => (x"87",x"ec",x"c1",x"c1"),
  1076 => (x"71",x"1e",x"4f",x"26"),
  1077 => (x"91",x"cb",x"49",x"4a"),
  1078 => (x"81",x"de",x"e4",x"c1"),
  1079 => (x"48",x"11",x"81",x"c8"),
  1080 => (x"58",x"c4",x"e8",x"c2"),
  1081 => (x"48",x"d8",x"e8",x"c2"),
  1082 => (x"49",x"c1",x"78",x"c0"),
  1083 => (x"26",x"87",x"df",x"dc"),
  1084 => (x"99",x"71",x"1e",x"4f"),
  1085 => (x"c1",x"87",x"d2",x"02"),
  1086 => (x"c0",x"48",x"f3",x"e5"),
  1087 => (x"c1",x"80",x"f7",x"50"),
  1088 => (x"c1",x"40",x"d2",x"c3"),
  1089 => (x"ce",x"78",x"d7",x"e4"),
  1090 => (x"ef",x"e5",x"c1",x"87"),
  1091 => (x"d0",x"e4",x"c1",x"48"),
  1092 => (x"c1",x"80",x"fc",x"78"),
  1093 => (x"26",x"78",x"c9",x"c3"),
  1094 => (x"5b",x"5e",x"0e",x"4f"),
  1095 => (x"f4",x"0e",x"5d",x"5c"),
  1096 => (x"ce",x"db",x"c2",x"86"),
  1097 => (x"c4",x"4c",x"c0",x"4d"),
  1098 => (x"78",x"c0",x"48",x"a6"),
  1099 => (x"bf",x"d8",x"e8",x"c2"),
  1100 => (x"06",x"a8",x"c0",x"48"),
  1101 => (x"c2",x"87",x"c0",x"c1"),
  1102 => (x"98",x"48",x"ce",x"db"),
  1103 => (x"87",x"f7",x"c0",x"02"),
  1104 => (x"1e",x"d3",x"f6",x"c0"),
  1105 => (x"c7",x"02",x"66",x"c8"),
  1106 => (x"48",x"a6",x"c4",x"87"),
  1107 => (x"87",x"c5",x"78",x"c0"),
  1108 => (x"c1",x"48",x"a6",x"c4"),
  1109 => (x"49",x"66",x"c4",x"78"),
  1110 => (x"c4",x"87",x"e6",x"e5"),
  1111 => (x"c1",x"4d",x"70",x"86"),
  1112 => (x"48",x"66",x"c4",x"84"),
  1113 => (x"a6",x"c8",x"80",x"c1"),
  1114 => (x"d8",x"e8",x"c2",x"58"),
  1115 => (x"c6",x"03",x"ac",x"bf"),
  1116 => (x"05",x"9d",x"75",x"87"),
  1117 => (x"c0",x"87",x"c9",x"ff"),
  1118 => (x"02",x"9d",x"75",x"4c"),
  1119 => (x"c0",x"87",x"dc",x"c3"),
  1120 => (x"c8",x"1e",x"d3",x"f6"),
  1121 => (x"87",x"c7",x"02",x"66"),
  1122 => (x"c0",x"48",x"a6",x"cc"),
  1123 => (x"cc",x"87",x"c5",x"78"),
  1124 => (x"78",x"c1",x"48",x"a6"),
  1125 => (x"e4",x"49",x"66",x"cc"),
  1126 => (x"86",x"c4",x"87",x"e7"),
  1127 => (x"98",x"48",x"7e",x"70"),
  1128 => (x"87",x"e4",x"c2",x"02"),
  1129 => (x"97",x"81",x"cb",x"49"),
  1130 => (x"99",x"d0",x"49",x"69"),
  1131 => (x"87",x"d4",x"c1",x"02"),
  1132 => (x"91",x"cb",x"49",x"74"),
  1133 => (x"81",x"de",x"e4",x"c1"),
  1134 => (x"79",x"e2",x"c2",x"c1"),
  1135 => (x"ff",x"c3",x"81",x"c8"),
  1136 => (x"de",x"49",x"74",x"51"),
  1137 => (x"ec",x"e8",x"c2",x"91"),
  1138 => (x"c2",x"85",x"71",x"4d"),
  1139 => (x"c1",x"7d",x"97",x"c1"),
  1140 => (x"e0",x"c0",x"49",x"a5"),
  1141 => (x"de",x"e3",x"c2",x"51"),
  1142 => (x"d2",x"02",x"bf",x"97"),
  1143 => (x"c2",x"84",x"c1",x"87"),
  1144 => (x"e3",x"c2",x"4b",x"a5"),
  1145 => (x"49",x"db",x"4a",x"de"),
  1146 => (x"87",x"fb",x"fa",x"fe"),
  1147 => (x"cd",x"87",x"d9",x"c1"),
  1148 => (x"51",x"c0",x"49",x"a5"),
  1149 => (x"a5",x"c2",x"84",x"c1"),
  1150 => (x"cb",x"4a",x"6e",x"4b"),
  1151 => (x"e6",x"fa",x"fe",x"49"),
  1152 => (x"87",x"c4",x"c1",x"87"),
  1153 => (x"91",x"cb",x"49",x"74"),
  1154 => (x"81",x"de",x"e4",x"c1"),
  1155 => (x"79",x"df",x"c0",x"c1"),
  1156 => (x"97",x"de",x"e3",x"c2"),
  1157 => (x"87",x"d8",x"02",x"bf"),
  1158 => (x"91",x"de",x"49",x"74"),
  1159 => (x"e8",x"c2",x"84",x"c1"),
  1160 => (x"83",x"71",x"4b",x"ec"),
  1161 => (x"4a",x"de",x"e3",x"c2"),
  1162 => (x"f9",x"fe",x"49",x"dd"),
  1163 => (x"87",x"d8",x"87",x"f9"),
  1164 => (x"93",x"de",x"4b",x"74"),
  1165 => (x"83",x"ec",x"e8",x"c2"),
  1166 => (x"c0",x"49",x"a3",x"cb"),
  1167 => (x"73",x"84",x"c1",x"51"),
  1168 => (x"49",x"cb",x"4a",x"6e"),
  1169 => (x"87",x"df",x"f9",x"fe"),
  1170 => (x"c1",x"48",x"66",x"c4"),
  1171 => (x"58",x"a6",x"c8",x"80"),
  1172 => (x"c0",x"03",x"ac",x"c7"),
  1173 => (x"05",x"6e",x"87",x"c5"),
  1174 => (x"74",x"87",x"e4",x"fc"),
  1175 => (x"f4",x"8e",x"f4",x"48"),
  1176 => (x"73",x"1e",x"87",x"f6"),
  1177 => (x"49",x"4b",x"71",x"1e"),
  1178 => (x"e4",x"c1",x"91",x"cb"),
  1179 => (x"a1",x"c8",x"81",x"de"),
  1180 => (x"ca",x"e4",x"c1",x"4a"),
  1181 => (x"c9",x"50",x"12",x"48"),
  1182 => (x"f9",x"c0",x"4a",x"a1"),
  1183 => (x"50",x"12",x"48",x"c0"),
  1184 => (x"e4",x"c1",x"81",x"ca"),
  1185 => (x"50",x"11",x"48",x"cb"),
  1186 => (x"97",x"cb",x"e4",x"c1"),
  1187 => (x"c0",x"1e",x"49",x"bf"),
  1188 => (x"87",x"cb",x"f5",x"49"),
  1189 => (x"48",x"c0",x"e8",x"c2"),
  1190 => (x"49",x"c1",x"78",x"de"),
  1191 => (x"26",x"87",x"ef",x"d5"),
  1192 => (x"0e",x"87",x"f9",x"f3"),
  1193 => (x"5d",x"5c",x"5b",x"5e"),
  1194 => (x"71",x"86",x"f4",x"0e"),
  1195 => (x"91",x"cb",x"49",x"4d"),
  1196 => (x"81",x"de",x"e4",x"c1"),
  1197 => (x"ca",x"4a",x"a1",x"c8"),
  1198 => (x"a6",x"c4",x"7e",x"a1"),
  1199 => (x"c8",x"ec",x"c2",x"48"),
  1200 => (x"97",x"6e",x"78",x"bf"),
  1201 => (x"66",x"c4",x"4b",x"bf"),
  1202 => (x"12",x"2c",x"73",x"4c"),
  1203 => (x"58",x"a6",x"cc",x"48"),
  1204 => (x"84",x"c1",x"9c",x"70"),
  1205 => (x"69",x"97",x"81",x"c9"),
  1206 => (x"04",x"ac",x"b7",x"49"),
  1207 => (x"4c",x"c0",x"87",x"c2"),
  1208 => (x"4a",x"bf",x"97",x"6e"),
  1209 => (x"72",x"49",x"66",x"c8"),
  1210 => (x"c4",x"b9",x"ff",x"31"),
  1211 => (x"48",x"74",x"99",x"66"),
  1212 => (x"4a",x"70",x"30",x"72"),
  1213 => (x"c2",x"b0",x"71",x"48"),
  1214 => (x"c0",x"58",x"cc",x"ec"),
  1215 => (x"c0",x"87",x"d8",x"e5"),
  1216 => (x"87",x"ca",x"d4",x"49"),
  1217 => (x"f7",x"c0",x"49",x"75"),
  1218 => (x"8e",x"f4",x"87",x"cd"),
  1219 => (x"1e",x"87",x"c9",x"f2"),
  1220 => (x"4b",x"71",x"1e",x"73"),
  1221 => (x"87",x"cb",x"fe",x"49"),
  1222 => (x"c6",x"fe",x"49",x"73"),
  1223 => (x"87",x"fc",x"f1",x"87"),
  1224 => (x"71",x"1e",x"73",x"1e"),
  1225 => (x"4a",x"a3",x"c6",x"4b"),
  1226 => (x"c1",x"87",x"db",x"02"),
  1227 => (x"87",x"d6",x"02",x"8a"),
  1228 => (x"da",x"c1",x"02",x"8a"),
  1229 => (x"c0",x"02",x"8a",x"87"),
  1230 => (x"02",x"8a",x"87",x"fc"),
  1231 => (x"8a",x"87",x"e1",x"c0"),
  1232 => (x"c1",x"87",x"cb",x"02"),
  1233 => (x"49",x"c7",x"87",x"db"),
  1234 => (x"c1",x"87",x"c7",x"f6"),
  1235 => (x"e8",x"c2",x"87",x"de"),
  1236 => (x"c1",x"02",x"bf",x"d8"),
  1237 => (x"c1",x"48",x"87",x"cb"),
  1238 => (x"dc",x"e8",x"c2",x"88"),
  1239 => (x"87",x"c1",x"c1",x"58"),
  1240 => (x"bf",x"dc",x"e8",x"c2"),
  1241 => (x"87",x"f9",x"c0",x"02"),
  1242 => (x"bf",x"d8",x"e8",x"c2"),
  1243 => (x"c2",x"80",x"c1",x"48"),
  1244 => (x"c0",x"58",x"dc",x"e8"),
  1245 => (x"e8",x"c2",x"87",x"eb"),
  1246 => (x"c6",x"49",x"bf",x"d8"),
  1247 => (x"dc",x"e8",x"c2",x"89"),
  1248 => (x"a9",x"b7",x"c0",x"59"),
  1249 => (x"c2",x"87",x"da",x"03"),
  1250 => (x"c0",x"48",x"d8",x"e8"),
  1251 => (x"c2",x"87",x"d2",x"78"),
  1252 => (x"02",x"bf",x"dc",x"e8"),
  1253 => (x"e8",x"c2",x"87",x"cb"),
  1254 => (x"c6",x"48",x"bf",x"d8"),
  1255 => (x"dc",x"e8",x"c2",x"80"),
  1256 => (x"d1",x"49",x"c0",x"58"),
  1257 => (x"49",x"73",x"87",x"e8"),
  1258 => (x"87",x"eb",x"f4",x"c0"),
  1259 => (x"0e",x"87",x"ed",x"ef"),
  1260 => (x"5d",x"5c",x"5b",x"5e"),
  1261 => (x"86",x"d4",x"ff",x"0e"),
  1262 => (x"c8",x"59",x"a6",x"dc"),
  1263 => (x"78",x"c0",x"48",x"a6"),
  1264 => (x"c0",x"c1",x"80",x"c4"),
  1265 => (x"80",x"c4",x"78",x"66"),
  1266 => (x"80",x"c4",x"78",x"c1"),
  1267 => (x"e8",x"c2",x"78",x"c1"),
  1268 => (x"78",x"c1",x"48",x"dc"),
  1269 => (x"bf",x"c0",x"e8",x"c2"),
  1270 => (x"05",x"a8",x"de",x"48"),
  1271 => (x"f8",x"f4",x"87",x"c9"),
  1272 => (x"58",x"a6",x"cc",x"87"),
  1273 => (x"e3",x"87",x"e6",x"cf"),
  1274 => (x"fb",x"e3",x"87",x"d9"),
  1275 => (x"87",x"c8",x"e3",x"87"),
  1276 => (x"fb",x"c0",x"4c",x"70"),
  1277 => (x"fb",x"c1",x"02",x"ac"),
  1278 => (x"05",x"66",x"d8",x"87"),
  1279 => (x"c0",x"87",x"ed",x"c1"),
  1280 => (x"c4",x"4a",x"66",x"fc"),
  1281 => (x"72",x"7e",x"6a",x"82"),
  1282 => (x"c2",x"e0",x"c1",x"1e"),
  1283 => (x"49",x"66",x"c4",x"48"),
  1284 => (x"20",x"4a",x"a1",x"c8"),
  1285 => (x"05",x"aa",x"71",x"41"),
  1286 => (x"51",x"10",x"87",x"f9"),
  1287 => (x"fc",x"c0",x"4a",x"26"),
  1288 => (x"c9",x"c1",x"48",x"66"),
  1289 => (x"49",x"6a",x"78",x"e2"),
  1290 => (x"51",x"74",x"81",x"c7"),
  1291 => (x"49",x"66",x"fc",x"c0"),
  1292 => (x"51",x"c1",x"81",x"c8"),
  1293 => (x"49",x"66",x"fc",x"c0"),
  1294 => (x"51",x"c0",x"81",x"c9"),
  1295 => (x"49",x"66",x"fc",x"c0"),
  1296 => (x"51",x"c0",x"81",x"ca"),
  1297 => (x"1e",x"d8",x"1e",x"c1"),
  1298 => (x"81",x"c8",x"49",x"6a"),
  1299 => (x"c8",x"87",x"ed",x"e2"),
  1300 => (x"66",x"c0",x"c1",x"86"),
  1301 => (x"01",x"a8",x"c0",x"48"),
  1302 => (x"a6",x"c8",x"87",x"c7"),
  1303 => (x"ce",x"78",x"c1",x"48"),
  1304 => (x"66",x"c0",x"c1",x"87"),
  1305 => (x"d0",x"88",x"c1",x"48"),
  1306 => (x"87",x"c3",x"58",x"a6"),
  1307 => (x"d0",x"87",x"f9",x"e1"),
  1308 => (x"78",x"c2",x"48",x"a6"),
  1309 => (x"cd",x"02",x"9c",x"74"),
  1310 => (x"66",x"c8",x"87",x"cf"),
  1311 => (x"66",x"c4",x"c1",x"48"),
  1312 => (x"c4",x"cd",x"03",x"a8"),
  1313 => (x"48",x"a6",x"dc",x"87"),
  1314 => (x"80",x"e8",x"78",x"c0"),
  1315 => (x"e7",x"e0",x"78",x"c0"),
  1316 => (x"c1",x"4c",x"70",x"87"),
  1317 => (x"c2",x"05",x"ac",x"d0"),
  1318 => (x"66",x"c4",x"87",x"d7"),
  1319 => (x"87",x"cb",x"e3",x"7e"),
  1320 => (x"e0",x"58",x"a6",x"c8"),
  1321 => (x"4c",x"70",x"87",x"d2"),
  1322 => (x"05",x"ac",x"ec",x"c0"),
  1323 => (x"c8",x"87",x"ed",x"c1"),
  1324 => (x"91",x"cb",x"49",x"66"),
  1325 => (x"81",x"66",x"fc",x"c0"),
  1326 => (x"6a",x"4a",x"a1",x"c4"),
  1327 => (x"4a",x"a1",x"c8",x"4d"),
  1328 => (x"c1",x"52",x"66",x"c4"),
  1329 => (x"ff",x"79",x"d2",x"c3"),
  1330 => (x"70",x"87",x"ed",x"df"),
  1331 => (x"d9",x"02",x"9c",x"4c"),
  1332 => (x"ac",x"fb",x"c0",x"87"),
  1333 => (x"74",x"87",x"d3",x"02"),
  1334 => (x"db",x"df",x"ff",x"55"),
  1335 => (x"9c",x"4c",x"70",x"87"),
  1336 => (x"c0",x"87",x"c7",x"02"),
  1337 => (x"ff",x"05",x"ac",x"fb"),
  1338 => (x"e0",x"c0",x"87",x"ed"),
  1339 => (x"55",x"c1",x"c2",x"55"),
  1340 => (x"d8",x"7d",x"97",x"c0"),
  1341 => (x"a8",x"6e",x"48",x"66"),
  1342 => (x"c8",x"87",x"db",x"05"),
  1343 => (x"66",x"cc",x"48",x"66"),
  1344 => (x"87",x"ca",x"04",x"a8"),
  1345 => (x"c1",x"48",x"66",x"c8"),
  1346 => (x"58",x"a6",x"cc",x"80"),
  1347 => (x"66",x"cc",x"87",x"c8"),
  1348 => (x"d0",x"88",x"c1",x"48"),
  1349 => (x"de",x"ff",x"58",x"a6"),
  1350 => (x"4c",x"70",x"87",x"de"),
  1351 => (x"05",x"ac",x"d0",x"c1"),
  1352 => (x"66",x"d4",x"87",x"c8"),
  1353 => (x"d8",x"80",x"c1",x"48"),
  1354 => (x"d0",x"c1",x"58",x"a6"),
  1355 => (x"e9",x"fd",x"02",x"ac"),
  1356 => (x"48",x"66",x"c4",x"87"),
  1357 => (x"05",x"a8",x"66",x"d8"),
  1358 => (x"c0",x"87",x"e0",x"c9"),
  1359 => (x"c0",x"48",x"a6",x"e0"),
  1360 => (x"c0",x"48",x"74",x"78"),
  1361 => (x"7e",x"70",x"88",x"fb"),
  1362 => (x"c9",x"02",x"98",x"48"),
  1363 => (x"cb",x"48",x"87",x"e2"),
  1364 => (x"48",x"7e",x"70",x"88"),
  1365 => (x"cd",x"c1",x"02",x"98"),
  1366 => (x"88",x"c9",x"48",x"87"),
  1367 => (x"98",x"48",x"7e",x"70"),
  1368 => (x"87",x"fe",x"c3",x"02"),
  1369 => (x"70",x"88",x"c4",x"48"),
  1370 => (x"02",x"98",x"48",x"7e"),
  1371 => (x"c1",x"48",x"87",x"ce"),
  1372 => (x"48",x"7e",x"70",x"88"),
  1373 => (x"e9",x"c3",x"02",x"98"),
  1374 => (x"87",x"d6",x"c8",x"87"),
  1375 => (x"c0",x"48",x"a6",x"dc"),
  1376 => (x"dc",x"ff",x"78",x"f0"),
  1377 => (x"4c",x"70",x"87",x"f2"),
  1378 => (x"02",x"ac",x"ec",x"c0"),
  1379 => (x"c0",x"87",x"c4",x"c0"),
  1380 => (x"c0",x"5c",x"a6",x"e0"),
  1381 => (x"cd",x"02",x"ac",x"ec"),
  1382 => (x"db",x"dc",x"ff",x"87"),
  1383 => (x"c0",x"4c",x"70",x"87"),
  1384 => (x"ff",x"05",x"ac",x"ec"),
  1385 => (x"ec",x"c0",x"87",x"f3"),
  1386 => (x"c4",x"c0",x"02",x"ac"),
  1387 => (x"c7",x"dc",x"ff",x"87"),
  1388 => (x"ca",x"1e",x"c0",x"87"),
  1389 => (x"49",x"66",x"d0",x"1e"),
  1390 => (x"c4",x"c1",x"91",x"cb"),
  1391 => (x"80",x"71",x"48",x"66"),
  1392 => (x"c8",x"58",x"a6",x"cc"),
  1393 => (x"80",x"c4",x"48",x"66"),
  1394 => (x"cc",x"58",x"a6",x"d0"),
  1395 => (x"ff",x"49",x"bf",x"66"),
  1396 => (x"c1",x"87",x"e9",x"dc"),
  1397 => (x"d4",x"1e",x"de",x"1e"),
  1398 => (x"ff",x"49",x"bf",x"66"),
  1399 => (x"d0",x"87",x"dd",x"dc"),
  1400 => (x"48",x"49",x"70",x"86"),
  1401 => (x"c0",x"88",x"08",x"c0"),
  1402 => (x"c0",x"58",x"a6",x"e8"),
  1403 => (x"ee",x"c0",x"06",x"a8"),
  1404 => (x"66",x"e4",x"c0",x"87"),
  1405 => (x"03",x"a8",x"dd",x"48"),
  1406 => (x"c4",x"87",x"e4",x"c0"),
  1407 => (x"c0",x"49",x"bf",x"66"),
  1408 => (x"c0",x"81",x"66",x"e4"),
  1409 => (x"e4",x"c0",x"51",x"e0"),
  1410 => (x"81",x"c1",x"49",x"66"),
  1411 => (x"81",x"bf",x"66",x"c4"),
  1412 => (x"c0",x"51",x"c1",x"c2"),
  1413 => (x"c2",x"49",x"66",x"e4"),
  1414 => (x"bf",x"66",x"c4",x"81"),
  1415 => (x"6e",x"51",x"c0",x"81"),
  1416 => (x"e2",x"c9",x"c1",x"48"),
  1417 => (x"c8",x"49",x"6e",x"78"),
  1418 => (x"51",x"66",x"d0",x"81"),
  1419 => (x"81",x"c9",x"49",x"6e"),
  1420 => (x"6e",x"51",x"66",x"d4"),
  1421 => (x"dc",x"81",x"ca",x"49"),
  1422 => (x"66",x"d0",x"51",x"66"),
  1423 => (x"d4",x"80",x"c1",x"48"),
  1424 => (x"66",x"c8",x"58",x"a6"),
  1425 => (x"a8",x"66",x"cc",x"48"),
  1426 => (x"87",x"cb",x"c0",x"04"),
  1427 => (x"c1",x"48",x"66",x"c8"),
  1428 => (x"58",x"a6",x"cc",x"80"),
  1429 => (x"cc",x"87",x"d9",x"c5"),
  1430 => (x"88",x"c1",x"48",x"66"),
  1431 => (x"c5",x"58",x"a6",x"d0"),
  1432 => (x"dc",x"ff",x"87",x"ce"),
  1433 => (x"e8",x"c0",x"87",x"c5"),
  1434 => (x"db",x"ff",x"58",x"a6"),
  1435 => (x"e0",x"c0",x"87",x"fd"),
  1436 => (x"ec",x"c0",x"58",x"a6"),
  1437 => (x"ca",x"c0",x"05",x"a8"),
  1438 => (x"48",x"a6",x"dc",x"87"),
  1439 => (x"78",x"66",x"e4",x"c0"),
  1440 => (x"ff",x"87",x"c4",x"c0"),
  1441 => (x"c8",x"87",x"f1",x"d8"),
  1442 => (x"91",x"cb",x"49",x"66"),
  1443 => (x"48",x"66",x"fc",x"c0"),
  1444 => (x"7e",x"70",x"80",x"71"),
  1445 => (x"6e",x"82",x"c8",x"4a"),
  1446 => (x"c0",x"81",x"ca",x"49"),
  1447 => (x"dc",x"51",x"66",x"e4"),
  1448 => (x"81",x"c1",x"49",x"66"),
  1449 => (x"89",x"66",x"e4",x"c0"),
  1450 => (x"30",x"71",x"48",x"c1"),
  1451 => (x"89",x"c1",x"49",x"70"),
  1452 => (x"c2",x"7a",x"97",x"71"),
  1453 => (x"49",x"bf",x"c8",x"ec"),
  1454 => (x"29",x"66",x"e4",x"c0"),
  1455 => (x"48",x"4a",x"6a",x"97"),
  1456 => (x"ec",x"c0",x"98",x"71"),
  1457 => (x"49",x"6e",x"58",x"a6"),
  1458 => (x"4d",x"69",x"81",x"c4"),
  1459 => (x"c4",x"48",x"66",x"d8"),
  1460 => (x"c0",x"02",x"a8",x"66"),
  1461 => (x"a6",x"c4",x"87",x"c8"),
  1462 => (x"c0",x"78",x"c0",x"48"),
  1463 => (x"a6",x"c4",x"87",x"c5"),
  1464 => (x"c4",x"78",x"c1",x"48"),
  1465 => (x"e0",x"c0",x"1e",x"66"),
  1466 => (x"ff",x"49",x"75",x"1e"),
  1467 => (x"c8",x"87",x"cd",x"d8"),
  1468 => (x"c0",x"4c",x"70",x"86"),
  1469 => (x"c1",x"06",x"ac",x"b7"),
  1470 => (x"85",x"74",x"87",x"d4"),
  1471 => (x"74",x"49",x"e0",x"c0"),
  1472 => (x"c1",x"4b",x"75",x"89"),
  1473 => (x"71",x"4a",x"cb",x"e0"),
  1474 => (x"87",x"db",x"e6",x"fe"),
  1475 => (x"e0",x"c0",x"85",x"c2"),
  1476 => (x"80",x"c1",x"48",x"66"),
  1477 => (x"58",x"a6",x"e4",x"c0"),
  1478 => (x"49",x"66",x"e8",x"c0"),
  1479 => (x"a9",x"70",x"81",x"c1"),
  1480 => (x"87",x"c8",x"c0",x"02"),
  1481 => (x"c0",x"48",x"a6",x"c4"),
  1482 => (x"87",x"c5",x"c0",x"78"),
  1483 => (x"c1",x"48",x"a6",x"c4"),
  1484 => (x"1e",x"66",x"c4",x"78"),
  1485 => (x"c0",x"49",x"a4",x"c2"),
  1486 => (x"88",x"71",x"48",x"e0"),
  1487 => (x"75",x"1e",x"49",x"70"),
  1488 => (x"f7",x"d6",x"ff",x"49"),
  1489 => (x"c0",x"86",x"c8",x"87"),
  1490 => (x"ff",x"01",x"a8",x"b7"),
  1491 => (x"e0",x"c0",x"87",x"c0"),
  1492 => (x"d1",x"c0",x"02",x"66"),
  1493 => (x"c9",x"49",x"6e",x"87"),
  1494 => (x"66",x"e0",x"c0",x"81"),
  1495 => (x"c1",x"48",x"6e",x"51"),
  1496 => (x"c0",x"78",x"e3",x"ca"),
  1497 => (x"49",x"6e",x"87",x"cc"),
  1498 => (x"51",x"c2",x"81",x"c9"),
  1499 => (x"cc",x"c1",x"48",x"6e"),
  1500 => (x"66",x"c8",x"78",x"cf"),
  1501 => (x"a8",x"66",x"cc",x"48"),
  1502 => (x"87",x"cb",x"c0",x"04"),
  1503 => (x"c1",x"48",x"66",x"c8"),
  1504 => (x"58",x"a6",x"cc",x"80"),
  1505 => (x"cc",x"87",x"e9",x"c0"),
  1506 => (x"88",x"c1",x"48",x"66"),
  1507 => (x"c0",x"58",x"a6",x"d0"),
  1508 => (x"d5",x"ff",x"87",x"de"),
  1509 => (x"4c",x"70",x"87",x"d2"),
  1510 => (x"c1",x"87",x"d5",x"c0"),
  1511 => (x"c0",x"05",x"ac",x"c6"),
  1512 => (x"66",x"d0",x"87",x"c8"),
  1513 => (x"d4",x"80",x"c1",x"48"),
  1514 => (x"d4",x"ff",x"58",x"a6"),
  1515 => (x"4c",x"70",x"87",x"fa"),
  1516 => (x"c1",x"48",x"66",x"d4"),
  1517 => (x"58",x"a6",x"d8",x"80"),
  1518 => (x"c0",x"02",x"9c",x"74"),
  1519 => (x"66",x"c8",x"87",x"cb"),
  1520 => (x"66",x"c4",x"c1",x"48"),
  1521 => (x"fc",x"f2",x"04",x"a8"),
  1522 => (x"d2",x"d4",x"ff",x"87"),
  1523 => (x"48",x"66",x"c8",x"87"),
  1524 => (x"c0",x"03",x"a8",x"c7"),
  1525 => (x"e8",x"c2",x"87",x"e5"),
  1526 => (x"78",x"c0",x"48",x"dc"),
  1527 => (x"cb",x"49",x"66",x"c8"),
  1528 => (x"66",x"fc",x"c0",x"91"),
  1529 => (x"4a",x"a1",x"c4",x"81"),
  1530 => (x"52",x"c0",x"4a",x"6a"),
  1531 => (x"48",x"66",x"c8",x"79"),
  1532 => (x"a6",x"cc",x"80",x"c1"),
  1533 => (x"04",x"a8",x"c7",x"58"),
  1534 => (x"ff",x"87",x"db",x"ff"),
  1535 => (x"de",x"ff",x"8e",x"d4"),
  1536 => (x"6f",x"4c",x"87",x"d6"),
  1537 => (x"2a",x"20",x"64",x"61"),
  1538 => (x"3a",x"00",x"20",x"2e"),
  1539 => (x"73",x"1e",x"00",x"20"),
  1540 => (x"9b",x"4b",x"71",x"1e"),
  1541 => (x"c2",x"87",x"c6",x"02"),
  1542 => (x"c0",x"48",x"d8",x"e8"),
  1543 => (x"c2",x"1e",x"c7",x"78"),
  1544 => (x"1e",x"bf",x"d8",x"e8"),
  1545 => (x"1e",x"de",x"e4",x"c1"),
  1546 => (x"bf",x"c0",x"e8",x"c2"),
  1547 => (x"87",x"ff",x"ed",x"49"),
  1548 => (x"e8",x"c2",x"86",x"cc"),
  1549 => (x"e2",x"49",x"bf",x"c0"),
  1550 => (x"9b",x"73",x"87",x"f7"),
  1551 => (x"c1",x"87",x"c8",x"02"),
  1552 => (x"c0",x"49",x"de",x"e4"),
  1553 => (x"ff",x"87",x"e2",x"e3"),
  1554 => (x"1e",x"87",x"d1",x"dd"),
  1555 => (x"4b",x"c0",x"1e",x"73"),
  1556 => (x"48",x"ca",x"e4",x"c1"),
  1557 => (x"e6",x"c1",x"50",x"c0"),
  1558 => (x"ff",x"49",x"bf",x"c1"),
  1559 => (x"70",x"87",x"e2",x"d7"),
  1560 => (x"87",x"c4",x"05",x"98"),
  1561 => (x"4b",x"ee",x"e1",x"c1"),
  1562 => (x"dc",x"ff",x"48",x"73"),
  1563 => (x"4f",x"52",x"87",x"ee"),
  1564 => (x"6f",x"6c",x"20",x"4d"),
  1565 => (x"6e",x"69",x"64",x"61"),
  1566 => (x"61",x"66",x"20",x"67"),
  1567 => (x"64",x"65",x"6c",x"69"),
  1568 => (x"e3",x"c7",x"1e",x"00"),
  1569 => (x"fe",x"49",x"c1",x"87"),
  1570 => (x"e9",x"fe",x"87",x"c4"),
  1571 => (x"98",x"70",x"87",x"c9"),
  1572 => (x"fe",x"87",x"cd",x"02"),
  1573 => (x"70",x"87",x"c3",x"f2"),
  1574 => (x"87",x"c4",x"02",x"98"),
  1575 => (x"87",x"c2",x"4a",x"c1"),
  1576 => (x"9a",x"72",x"4a",x"c0"),
  1577 => (x"c0",x"87",x"ce",x"05"),
  1578 => (x"d1",x"e3",x"c1",x"1e"),
  1579 => (x"ee",x"ee",x"c0",x"49"),
  1580 => (x"fe",x"86",x"c4",x"87"),
  1581 => (x"c1",x"1e",x"c0",x"87"),
  1582 => (x"c0",x"49",x"dc",x"e3"),
  1583 => (x"c0",x"87",x"e0",x"ee"),
  1584 => (x"87",x"c7",x"fe",x"1e"),
  1585 => (x"ee",x"c0",x"49",x"70"),
  1586 => (x"da",x"c3",x"87",x"d5"),
  1587 => (x"26",x"8e",x"f8",x"87"),
  1588 => (x"20",x"44",x"53",x"4f"),
  1589 => (x"6c",x"69",x"61",x"66"),
  1590 => (x"00",x"2e",x"64",x"65"),
  1591 => (x"74",x"6f",x"6f",x"42"),
  1592 => (x"2e",x"67",x"6e",x"69"),
  1593 => (x"1e",x"00",x"2e",x"2e"),
  1594 => (x"87",x"fa",x"e5",x"c0"),
  1595 => (x"87",x"e9",x"f1",x"c0"),
  1596 => (x"4f",x"26",x"87",x"f6"),
  1597 => (x"d8",x"e8",x"c2",x"1e"),
  1598 => (x"c2",x"78",x"c0",x"48"),
  1599 => (x"c0",x"48",x"c0",x"e8"),
  1600 => (x"87",x"fd",x"fd",x"78"),
  1601 => (x"48",x"c0",x"87",x"e1"),
  1602 => (x"00",x"00",x"4f",x"26"),
  1603 => (x"00",x"00",x"00",x"01"),
  1604 => (x"78",x"45",x"20",x"80"),
  1605 => (x"80",x"00",x"74",x"69"),
  1606 => (x"63",x"61",x"42",x"20"),
  1607 => (x"10",x"1f",x"00",x"6b"),
  1608 => (x"2a",x"2c",x"00",x"00"),
  1609 => (x"00",x"00",x"00",x"00"),
  1610 => (x"00",x"10",x"1f",x"00"),
  1611 => (x"00",x"2a",x"4a",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"00",x"10",x"1f"),
  1614 => (x"00",x"00",x"2a",x"68"),
  1615 => (x"1f",x"00",x"00",x"00"),
  1616 => (x"86",x"00",x"00",x"10"),
  1617 => (x"00",x"00",x"00",x"2a"),
  1618 => (x"10",x"1f",x"00",x"00"),
  1619 => (x"2a",x"a4",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"10",x"1f",x"00"),
  1622 => (x"00",x"2a",x"c2",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"00",x"10",x"1f"),
  1625 => (x"00",x"00",x"2a",x"e0"),
  1626 => (x"d2",x"00",x"00",x"00"),
  1627 => (x"00",x"00",x"00",x"10"),
  1628 => (x"00",x"00",x"00",x"00"),
  1629 => (x"13",x"20",x"00",x"00"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"00",x"00",x"00",x"00"),
  1632 => (x"00",x"19",x"85",x"00"),
  1633 => (x"39",x"49",x"54",x"00"),
  1634 => (x"20",x"41",x"34",x"39"),
  1635 => (x"4d",x"4f",x"52",x"20"),
  1636 => (x"f0",x"fe",x"1e",x"00"),
  1637 => (x"cd",x"78",x"c0",x"48"),
  1638 => (x"26",x"09",x"79",x"09"),
  1639 => (x"fe",x"1e",x"1e",x"4f"),
  1640 => (x"48",x"7e",x"bf",x"f0"),
  1641 => (x"1e",x"4f",x"26",x"26"),
  1642 => (x"c1",x"48",x"f0",x"fe"),
  1643 => (x"1e",x"4f",x"26",x"78"),
  1644 => (x"c0",x"48",x"f0",x"fe"),
  1645 => (x"1e",x"4f",x"26",x"78"),
  1646 => (x"52",x"c0",x"4a",x"71"),
  1647 => (x"0e",x"4f",x"26",x"52"),
  1648 => (x"5d",x"5c",x"5b",x"5e"),
  1649 => (x"71",x"86",x"f4",x"0e"),
  1650 => (x"7e",x"6d",x"97",x"4d"),
  1651 => (x"97",x"4c",x"a5",x"c1"),
  1652 => (x"a6",x"c8",x"48",x"6c"),
  1653 => (x"c4",x"48",x"6e",x"58"),
  1654 => (x"c5",x"05",x"a8",x"66"),
  1655 => (x"c0",x"48",x"ff",x"87"),
  1656 => (x"ca",x"ff",x"87",x"e6"),
  1657 => (x"49",x"a5",x"c2",x"87"),
  1658 => (x"71",x"4b",x"6c",x"97"),
  1659 => (x"6b",x"97",x"4b",x"a3"),
  1660 => (x"7e",x"6c",x"97",x"4b"),
  1661 => (x"80",x"c1",x"48",x"6e"),
  1662 => (x"c7",x"58",x"a6",x"c8"),
  1663 => (x"58",x"a6",x"cc",x"98"),
  1664 => (x"fe",x"7c",x"97",x"70"),
  1665 => (x"48",x"73",x"87",x"e1"),
  1666 => (x"4d",x"26",x"8e",x"f4"),
  1667 => (x"4b",x"26",x"4c",x"26"),
  1668 => (x"5e",x"0e",x"4f",x"26"),
  1669 => (x"f4",x"0e",x"5c",x"5b"),
  1670 => (x"d8",x"4c",x"71",x"86"),
  1671 => (x"ff",x"c3",x"4a",x"66"),
  1672 => (x"4b",x"a4",x"c2",x"9a"),
  1673 => (x"73",x"49",x"6c",x"97"),
  1674 => (x"51",x"72",x"49",x"a1"),
  1675 => (x"6e",x"7e",x"6c",x"97"),
  1676 => (x"c8",x"80",x"c1",x"48"),
  1677 => (x"98",x"c7",x"58",x"a6"),
  1678 => (x"70",x"58",x"a6",x"cc"),
  1679 => (x"ff",x"8e",x"f4",x"54"),
  1680 => (x"1e",x"1e",x"87",x"ca"),
  1681 => (x"e0",x"87",x"e8",x"fd"),
  1682 => (x"c0",x"49",x"4a",x"bf"),
  1683 => (x"02",x"99",x"c0",x"e0"),
  1684 => (x"1e",x"72",x"87",x"cb"),
  1685 => (x"49",x"fe",x"eb",x"c2"),
  1686 => (x"c4",x"87",x"f7",x"fe"),
  1687 => (x"87",x"fd",x"fc",x"86"),
  1688 => (x"c2",x"fd",x"7e",x"70"),
  1689 => (x"4f",x"26",x"26",x"87"),
  1690 => (x"fe",x"eb",x"c2",x"1e"),
  1691 => (x"87",x"c7",x"fd",x"49"),
  1692 => (x"49",x"c2",x"e9",x"c1"),
  1693 => (x"c3",x"87",x"da",x"fc"),
  1694 => (x"4f",x"26",x"87",x"f7"),
  1695 => (x"5c",x"5b",x"5e",x"0e"),
  1696 => (x"4d",x"71",x"0e",x"5d"),
  1697 => (x"49",x"fe",x"eb",x"c2"),
  1698 => (x"70",x"87",x"f4",x"fc"),
  1699 => (x"ab",x"b7",x"c0",x"4b"),
  1700 => (x"87",x"c2",x"c3",x"04"),
  1701 => (x"05",x"ab",x"f0",x"c3"),
  1702 => (x"ed",x"c1",x"87",x"c9"),
  1703 => (x"78",x"c1",x"48",x"e0"),
  1704 => (x"c3",x"87",x"e3",x"c2"),
  1705 => (x"c9",x"05",x"ab",x"e0"),
  1706 => (x"e4",x"ed",x"c1",x"87"),
  1707 => (x"c2",x"78",x"c1",x"48"),
  1708 => (x"ed",x"c1",x"87",x"d4"),
  1709 => (x"c6",x"02",x"bf",x"e4"),
  1710 => (x"a3",x"c0",x"c2",x"87"),
  1711 => (x"73",x"87",x"c2",x"4c"),
  1712 => (x"e0",x"ed",x"c1",x"4c"),
  1713 => (x"e0",x"c0",x"02",x"bf"),
  1714 => (x"c4",x"49",x"74",x"87"),
  1715 => (x"c1",x"91",x"29",x"b7"),
  1716 => (x"74",x"81",x"c0",x"ef"),
  1717 => (x"c2",x"9a",x"cf",x"4a"),
  1718 => (x"72",x"48",x"c1",x"92"),
  1719 => (x"ff",x"4a",x"70",x"30"),
  1720 => (x"69",x"48",x"72",x"ba"),
  1721 => (x"db",x"79",x"70",x"98"),
  1722 => (x"c4",x"49",x"74",x"87"),
  1723 => (x"c1",x"91",x"29",x"b7"),
  1724 => (x"74",x"81",x"c0",x"ef"),
  1725 => (x"c2",x"9a",x"cf",x"4a"),
  1726 => (x"72",x"48",x"c3",x"92"),
  1727 => (x"48",x"4a",x"70",x"30"),
  1728 => (x"79",x"70",x"b0",x"69"),
  1729 => (x"c0",x"05",x"9d",x"75"),
  1730 => (x"d0",x"ff",x"87",x"f0"),
  1731 => (x"78",x"e1",x"c8",x"48"),
  1732 => (x"c5",x"48",x"d4",x"ff"),
  1733 => (x"e4",x"ed",x"c1",x"78"),
  1734 => (x"87",x"c3",x"02",x"bf"),
  1735 => (x"c1",x"78",x"e0",x"c3"),
  1736 => (x"02",x"bf",x"e0",x"ed"),
  1737 => (x"d4",x"ff",x"87",x"c6"),
  1738 => (x"78",x"f0",x"c3",x"48"),
  1739 => (x"7b",x"0b",x"d4",x"ff"),
  1740 => (x"48",x"d0",x"ff",x"0b"),
  1741 => (x"c0",x"78",x"e1",x"c8"),
  1742 => (x"ed",x"c1",x"78",x"e0"),
  1743 => (x"78",x"c0",x"48",x"e4"),
  1744 => (x"48",x"e0",x"ed",x"c1"),
  1745 => (x"eb",x"c2",x"78",x"c0"),
  1746 => (x"f2",x"f9",x"49",x"fe"),
  1747 => (x"c0",x"4b",x"70",x"87"),
  1748 => (x"fc",x"03",x"ab",x"b7"),
  1749 => (x"48",x"c0",x"87",x"fe"),
  1750 => (x"4c",x"26",x"4d",x"26"),
  1751 => (x"4f",x"26",x"4b",x"26"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"49",x"4a",x"71",x"1e"),
  1755 => (x"26",x"87",x"cd",x"fc"),
  1756 => (x"4a",x"c0",x"1e",x"4f"),
  1757 => (x"91",x"c4",x"49",x"72"),
  1758 => (x"81",x"c0",x"ef",x"c1"),
  1759 => (x"82",x"c1",x"79",x"c0"),
  1760 => (x"04",x"aa",x"b7",x"d0"),
  1761 => (x"4f",x"26",x"87",x"ee"),
  1762 => (x"5c",x"5b",x"5e",x"0e"),
  1763 => (x"4d",x"71",x"0e",x"5d"),
  1764 => (x"75",x"87",x"dc",x"f8"),
  1765 => (x"2a",x"b7",x"c4",x"4a"),
  1766 => (x"c0",x"ef",x"c1",x"92"),
  1767 => (x"cf",x"4c",x"75",x"82"),
  1768 => (x"6a",x"94",x"c2",x"9c"),
  1769 => (x"2b",x"74",x"4b",x"49"),
  1770 => (x"48",x"c2",x"9b",x"c3"),
  1771 => (x"4c",x"70",x"30",x"74"),
  1772 => (x"48",x"74",x"bc",x"ff"),
  1773 => (x"7a",x"70",x"98",x"71"),
  1774 => (x"73",x"87",x"ec",x"f7"),
  1775 => (x"87",x"d8",x"fe",x"48"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"48",x"d0",x"ff",x"1e"),
  1793 => (x"71",x"78",x"e1",x"c8"),
  1794 => (x"08",x"d4",x"ff",x"48"),
  1795 => (x"1e",x"4f",x"26",x"78"),
  1796 => (x"c8",x"48",x"d0",x"ff"),
  1797 => (x"48",x"71",x"78",x"e1"),
  1798 => (x"78",x"08",x"d4",x"ff"),
  1799 => (x"ff",x"48",x"66",x"c4"),
  1800 => (x"26",x"78",x"08",x"d4"),
  1801 => (x"4a",x"71",x"1e",x"4f"),
  1802 => (x"1e",x"49",x"66",x"c4"),
  1803 => (x"de",x"ff",x"49",x"72"),
  1804 => (x"48",x"d0",x"ff",x"87"),
  1805 => (x"26",x"78",x"e0",x"c0"),
  1806 => (x"73",x"1e",x"4f",x"26"),
  1807 => (x"c8",x"4b",x"71",x"1e"),
  1808 => (x"73",x"1e",x"49",x"66"),
  1809 => (x"a2",x"e0",x"c1",x"4a"),
  1810 => (x"87",x"d9",x"ff",x"49"),
  1811 => (x"26",x"87",x"c4",x"26"),
  1812 => (x"26",x"4c",x"26",x"4d"),
  1813 => (x"1e",x"4f",x"26",x"4b"),
  1814 => (x"c3",x"4a",x"d4",x"ff"),
  1815 => (x"d0",x"ff",x"7a",x"ff"),
  1816 => (x"78",x"e1",x"c0",x"48"),
  1817 => (x"ec",x"c2",x"7a",x"de"),
  1818 => (x"49",x"7a",x"bf",x"c8"),
  1819 => (x"70",x"28",x"c8",x"48"),
  1820 => (x"d0",x"48",x"71",x"7a"),
  1821 => (x"71",x"7a",x"70",x"28"),
  1822 => (x"70",x"28",x"d8",x"48"),
  1823 => (x"48",x"d0",x"ff",x"7a"),
  1824 => (x"26",x"78",x"e0",x"c0"),
  1825 => (x"d0",x"ff",x"1e",x"4f"),
  1826 => (x"78",x"c9",x"c8",x"48"),
  1827 => (x"d4",x"ff",x"48",x"71"),
  1828 => (x"4f",x"26",x"78",x"08"),
  1829 => (x"49",x"4a",x"71",x"1e"),
  1830 => (x"d0",x"ff",x"87",x"eb"),
  1831 => (x"26",x"78",x"c8",x"48"),
  1832 => (x"1e",x"73",x"1e",x"4f"),
  1833 => (x"ec",x"c2",x"4b",x"71"),
  1834 => (x"c3",x"02",x"bf",x"d8"),
  1835 => (x"87",x"eb",x"c2",x"87"),
  1836 => (x"c8",x"48",x"d0",x"ff"),
  1837 => (x"48",x"73",x"78",x"c9"),
  1838 => (x"ff",x"b0",x"e0",x"c0"),
  1839 => (x"c2",x"78",x"08",x"d4"),
  1840 => (x"c0",x"48",x"cc",x"ec"),
  1841 => (x"02",x"66",x"c8",x"78"),
  1842 => (x"ff",x"c3",x"87",x"c5"),
  1843 => (x"c0",x"87",x"c2",x"49"),
  1844 => (x"d4",x"ec",x"c2",x"49"),
  1845 => (x"02",x"66",x"cc",x"59"),
  1846 => (x"d5",x"c5",x"87",x"c6"),
  1847 => (x"87",x"c4",x"4a",x"d5"),
  1848 => (x"4a",x"ff",x"ff",x"cf"),
  1849 => (x"5a",x"d8",x"ec",x"c2"),
  1850 => (x"48",x"d8",x"ec",x"c2"),
  1851 => (x"87",x"c4",x"78",x"c1"),
  1852 => (x"4c",x"26",x"4d",x"26"),
  1853 => (x"4f",x"26",x"4b",x"26"),
  1854 => (x"5c",x"5b",x"5e",x"0e"),
  1855 => (x"4a",x"71",x"0e",x"5d"),
  1856 => (x"bf",x"d4",x"ec",x"c2"),
  1857 => (x"02",x"9a",x"72",x"4c"),
  1858 => (x"c8",x"49",x"87",x"cb"),
  1859 => (x"d7",x"f2",x"c1",x"91"),
  1860 => (x"c4",x"83",x"71",x"4b"),
  1861 => (x"d7",x"f6",x"c1",x"87"),
  1862 => (x"13",x"4d",x"c0",x"4b"),
  1863 => (x"c2",x"99",x"74",x"49"),
  1864 => (x"48",x"bf",x"d0",x"ec"),
  1865 => (x"d4",x"ff",x"b8",x"71"),
  1866 => (x"b7",x"c1",x"78",x"08"),
  1867 => (x"b7",x"c8",x"85",x"2c"),
  1868 => (x"87",x"e7",x"04",x"ad"),
  1869 => (x"bf",x"cc",x"ec",x"c2"),
  1870 => (x"c2",x"80",x"c8",x"48"),
  1871 => (x"fe",x"58",x"d0",x"ec"),
  1872 => (x"73",x"1e",x"87",x"ee"),
  1873 => (x"13",x"4b",x"71",x"1e"),
  1874 => (x"cb",x"02",x"9a",x"4a"),
  1875 => (x"fe",x"49",x"72",x"87"),
  1876 => (x"4a",x"13",x"87",x"e6"),
  1877 => (x"87",x"f5",x"05",x"9a"),
  1878 => (x"1e",x"87",x"d9",x"fe"),
  1879 => (x"bf",x"cc",x"ec",x"c2"),
  1880 => (x"cc",x"ec",x"c2",x"49"),
  1881 => (x"78",x"a1",x"c1",x"48"),
  1882 => (x"a9",x"b7",x"c0",x"c4"),
  1883 => (x"ff",x"87",x"db",x"03"),
  1884 => (x"ec",x"c2",x"48",x"d4"),
  1885 => (x"c2",x"78",x"bf",x"d0"),
  1886 => (x"49",x"bf",x"cc",x"ec"),
  1887 => (x"48",x"cc",x"ec",x"c2"),
  1888 => (x"c4",x"78",x"a1",x"c1"),
  1889 => (x"04",x"a9",x"b7",x"c0"),
  1890 => (x"d0",x"ff",x"87",x"e5"),
  1891 => (x"c2",x"78",x"c8",x"48"),
  1892 => (x"c0",x"48",x"d8",x"ec"),
  1893 => (x"00",x"4f",x"26",x"78"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"5f",x"5f",x"00",x"00"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"03",x"00",x"03",x"03"),
  1899 => (x"14",x"00",x"00",x"03"),
  1900 => (x"7f",x"14",x"7f",x"7f"),
  1901 => (x"00",x"00",x"14",x"7f"),
  1902 => (x"6b",x"6b",x"2e",x"24"),
  1903 => (x"4c",x"00",x"12",x"3a"),
  1904 => (x"6c",x"18",x"36",x"6a"),
  1905 => (x"30",x"00",x"32",x"56"),
  1906 => (x"77",x"59",x"4f",x"7e"),
  1907 => (x"00",x"40",x"68",x"3a"),
  1908 => (x"03",x"07",x"04",x"00"),
  1909 => (x"00",x"00",x"00",x"00"),
  1910 => (x"63",x"3e",x"1c",x"00"),
  1911 => (x"00",x"00",x"00",x"41"),
  1912 => (x"3e",x"63",x"41",x"00"),
  1913 => (x"08",x"00",x"00",x"1c"),
  1914 => (x"1c",x"1c",x"3e",x"2a"),
  1915 => (x"00",x"08",x"2a",x"3e"),
  1916 => (x"3e",x"3e",x"08",x"08"),
  1917 => (x"00",x"00",x"08",x"08"),
  1918 => (x"60",x"e0",x"80",x"00"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"08",x"08",x"08",x"08"),
  1921 => (x"00",x"00",x"08",x"08"),
  1922 => (x"60",x"60",x"00",x"00"),
  1923 => (x"40",x"00",x"00",x"00"),
  1924 => (x"0c",x"18",x"30",x"60"),
  1925 => (x"00",x"01",x"03",x"06"),
  1926 => (x"4d",x"59",x"7f",x"3e"),
  1927 => (x"00",x"00",x"3e",x"7f"),
  1928 => (x"7f",x"7f",x"06",x"04"),
  1929 => (x"00",x"00",x"00",x"00"),
  1930 => (x"59",x"71",x"63",x"42"),
  1931 => (x"00",x"00",x"46",x"4f"),
  1932 => (x"49",x"49",x"63",x"22"),
  1933 => (x"18",x"00",x"36",x"7f"),
  1934 => (x"7f",x"13",x"16",x"1c"),
  1935 => (x"00",x"00",x"10",x"7f"),
  1936 => (x"45",x"45",x"67",x"27"),
  1937 => (x"00",x"00",x"39",x"7d"),
  1938 => (x"49",x"4b",x"7e",x"3c"),
  1939 => (x"00",x"00",x"30",x"79"),
  1940 => (x"79",x"71",x"01",x"01"),
  1941 => (x"00",x"00",x"07",x"0f"),
  1942 => (x"49",x"49",x"7f",x"36"),
  1943 => (x"00",x"00",x"36",x"7f"),
  1944 => (x"69",x"49",x"4f",x"06"),
  1945 => (x"00",x"00",x"1e",x"3f"),
  1946 => (x"66",x"66",x"00",x"00"),
  1947 => (x"00",x"00",x"00",x"00"),
  1948 => (x"66",x"e6",x"80",x"00"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"14",x"14",x"08",x"08"),
  1951 => (x"00",x"00",x"22",x"22"),
  1952 => (x"14",x"14",x"14",x"14"),
  1953 => (x"00",x"00",x"14",x"14"),
  1954 => (x"14",x"14",x"22",x"22"),
  1955 => (x"00",x"00",x"08",x"08"),
  1956 => (x"59",x"51",x"03",x"02"),
  1957 => (x"3e",x"00",x"06",x"0f"),
  1958 => (x"55",x"5d",x"41",x"7f"),
  1959 => (x"00",x"00",x"1e",x"1f"),
  1960 => (x"09",x"09",x"7f",x"7e"),
  1961 => (x"00",x"00",x"7e",x"7f"),
  1962 => (x"49",x"49",x"7f",x"7f"),
  1963 => (x"00",x"00",x"36",x"7f"),
  1964 => (x"41",x"63",x"3e",x"1c"),
  1965 => (x"00",x"00",x"41",x"41"),
  1966 => (x"63",x"41",x"7f",x"7f"),
  1967 => (x"00",x"00",x"1c",x"3e"),
  1968 => (x"49",x"49",x"7f",x"7f"),
  1969 => (x"00",x"00",x"41",x"41"),
  1970 => (x"09",x"09",x"7f",x"7f"),
  1971 => (x"00",x"00",x"01",x"01"),
  1972 => (x"49",x"41",x"7f",x"3e"),
  1973 => (x"00",x"00",x"7a",x"7b"),
  1974 => (x"08",x"08",x"7f",x"7f"),
  1975 => (x"00",x"00",x"7f",x"7f"),
  1976 => (x"7f",x"7f",x"41",x"00"),
  1977 => (x"00",x"00",x"00",x"41"),
  1978 => (x"40",x"40",x"60",x"20"),
  1979 => (x"7f",x"00",x"3f",x"7f"),
  1980 => (x"36",x"1c",x"08",x"7f"),
  1981 => (x"00",x"00",x"41",x"63"),
  1982 => (x"40",x"40",x"7f",x"7f"),
  1983 => (x"7f",x"00",x"40",x"40"),
  1984 => (x"06",x"0c",x"06",x"7f"),
  1985 => (x"7f",x"00",x"7f",x"7f"),
  1986 => (x"18",x"0c",x"06",x"7f"),
  1987 => (x"00",x"00",x"7f",x"7f"),
  1988 => (x"41",x"41",x"7f",x"3e"),
  1989 => (x"00",x"00",x"3e",x"7f"),
  1990 => (x"09",x"09",x"7f",x"7f"),
  1991 => (x"3e",x"00",x"06",x"0f"),
  1992 => (x"7f",x"61",x"41",x"7f"),
  1993 => (x"00",x"00",x"40",x"7e"),
  1994 => (x"19",x"09",x"7f",x"7f"),
  1995 => (x"00",x"00",x"66",x"7f"),
  1996 => (x"59",x"4d",x"6f",x"26"),
  1997 => (x"00",x"00",x"32",x"7b"),
  1998 => (x"7f",x"7f",x"01",x"01"),
  1999 => (x"00",x"00",x"01",x"01"),
  2000 => (x"40",x"40",x"7f",x"3f"),
  2001 => (x"00",x"00",x"3f",x"7f"),
  2002 => (x"70",x"70",x"3f",x"0f"),
  2003 => (x"7f",x"00",x"0f",x"3f"),
  2004 => (x"30",x"18",x"30",x"7f"),
  2005 => (x"41",x"00",x"7f",x"7f"),
  2006 => (x"1c",x"1c",x"36",x"63"),
  2007 => (x"01",x"41",x"63",x"36"),
  2008 => (x"7c",x"7c",x"06",x"03"),
  2009 => (x"61",x"01",x"03",x"06"),
  2010 => (x"47",x"4d",x"59",x"71"),
  2011 => (x"00",x"00",x"41",x"43"),
  2012 => (x"41",x"7f",x"7f",x"00"),
  2013 => (x"01",x"00",x"00",x"41"),
  2014 => (x"18",x"0c",x"06",x"03"),
  2015 => (x"00",x"40",x"60",x"30"),
  2016 => (x"7f",x"41",x"41",x"00"),
  2017 => (x"08",x"00",x"00",x"7f"),
  2018 => (x"06",x"03",x"06",x"0c"),
  2019 => (x"80",x"00",x"08",x"0c"),
  2020 => (x"80",x"80",x"80",x"80"),
  2021 => (x"00",x"00",x"80",x"80"),
  2022 => (x"07",x"03",x"00",x"00"),
  2023 => (x"00",x"00",x"00",x"04"),
  2024 => (x"54",x"54",x"74",x"20"),
  2025 => (x"00",x"00",x"78",x"7c"),
  2026 => (x"44",x"44",x"7f",x"7f"),
  2027 => (x"00",x"00",x"38",x"7c"),
  2028 => (x"44",x"44",x"7c",x"38"),
  2029 => (x"00",x"00",x"00",x"44"),
  2030 => (x"44",x"44",x"7c",x"38"),
  2031 => (x"00",x"00",x"7f",x"7f"),
  2032 => (x"54",x"54",x"7c",x"38"),
  2033 => (x"00",x"00",x"18",x"5c"),
  2034 => (x"05",x"7f",x"7e",x"04"),
  2035 => (x"00",x"00",x"00",x"05"),
  2036 => (x"a4",x"a4",x"bc",x"18"),
  2037 => (x"00",x"00",x"7c",x"fc"),
  2038 => (x"04",x"04",x"7f",x"7f"),
  2039 => (x"00",x"00",x"78",x"7c"),
  2040 => (x"7d",x"3d",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"40"),
  2042 => (x"fd",x"80",x"80",x"80"),
  2043 => (x"00",x"00",x"00",x"7d"),
  2044 => (x"38",x"10",x"7f",x"7f"),
  2045 => (x"00",x"00",x"44",x"6c"),
  2046 => (x"7f",x"3f",x"00",x"00"),
  2047 => (x"7c",x"00",x"00",x"40"),
  2048 => (x"0c",x"18",x"0c",x"7c"),
  2049 => (x"00",x"00",x"78",x"7c"),
  2050 => (x"04",x"04",x"7c",x"7c"),
  2051 => (x"00",x"00",x"78",x"7c"),
  2052 => (x"44",x"44",x"7c",x"38"),
  2053 => (x"00",x"00",x"38",x"7c"),
  2054 => (x"24",x"24",x"fc",x"fc"),
  2055 => (x"00",x"00",x"18",x"3c"),
  2056 => (x"24",x"24",x"3c",x"18"),
  2057 => (x"00",x"00",x"fc",x"fc"),
  2058 => (x"04",x"04",x"7c",x"7c"),
  2059 => (x"00",x"00",x"08",x"0c"),
  2060 => (x"54",x"54",x"5c",x"48"),
  2061 => (x"00",x"00",x"20",x"74"),
  2062 => (x"44",x"7f",x"3f",x"04"),
  2063 => (x"00",x"00",x"00",x"44"),
  2064 => (x"40",x"40",x"7c",x"3c"),
  2065 => (x"00",x"00",x"7c",x"7c"),
  2066 => (x"60",x"60",x"3c",x"1c"),
  2067 => (x"3c",x"00",x"1c",x"3c"),
  2068 => (x"60",x"30",x"60",x"7c"),
  2069 => (x"44",x"00",x"3c",x"7c"),
  2070 => (x"38",x"10",x"38",x"6c"),
  2071 => (x"00",x"00",x"44",x"6c"),
  2072 => (x"60",x"e0",x"bc",x"1c"),
  2073 => (x"00",x"00",x"1c",x"3c"),
  2074 => (x"5c",x"74",x"64",x"44"),
  2075 => (x"00",x"00",x"44",x"4c"),
  2076 => (x"77",x"3e",x"08",x"08"),
  2077 => (x"00",x"00",x"41",x"41"),
  2078 => (x"7f",x"7f",x"00",x"00"),
  2079 => (x"00",x"00",x"00",x"00"),
  2080 => (x"3e",x"77",x"41",x"41"),
  2081 => (x"02",x"00",x"08",x"08"),
  2082 => (x"02",x"03",x"01",x"01"),
  2083 => (x"7f",x"00",x"01",x"02"),
  2084 => (x"7f",x"7f",x"7f",x"7f"),
  2085 => (x"08",x"00",x"7f",x"7f"),
  2086 => (x"3e",x"1c",x"1c",x"08"),
  2087 => (x"7f",x"7f",x"7f",x"3e"),
  2088 => (x"1c",x"3e",x"3e",x"7f"),
  2089 => (x"00",x"08",x"08",x"1c"),
  2090 => (x"7c",x"7c",x"18",x"10"),
  2091 => (x"00",x"00",x"10",x"18"),
  2092 => (x"7c",x"7c",x"30",x"10"),
  2093 => (x"10",x"00",x"10",x"30"),
  2094 => (x"78",x"60",x"60",x"30"),
  2095 => (x"42",x"00",x"06",x"1e"),
  2096 => (x"3c",x"18",x"3c",x"66"),
  2097 => (x"78",x"00",x"42",x"66"),
  2098 => (x"c6",x"c2",x"6a",x"38"),
  2099 => (x"60",x"00",x"38",x"6c"),
  2100 => (x"00",x"60",x"00",x"00"),
  2101 => (x"0e",x"00",x"60",x"00"),
  2102 => (x"5d",x"5c",x"5b",x"5e"),
  2103 => (x"4c",x"71",x"1e",x"0e"),
  2104 => (x"bf",x"e9",x"ec",x"c2"),
  2105 => (x"c0",x"4b",x"c0",x"4d"),
  2106 => (x"02",x"ab",x"74",x"1e"),
  2107 => (x"a6",x"c4",x"87",x"c7"),
  2108 => (x"c5",x"78",x"c0",x"48"),
  2109 => (x"48",x"a6",x"c4",x"87"),
  2110 => (x"66",x"c4",x"78",x"c1"),
  2111 => (x"ee",x"49",x"73",x"1e"),
  2112 => (x"86",x"c8",x"87",x"df"),
  2113 => (x"ef",x"49",x"e0",x"c0"),
  2114 => (x"a5",x"c4",x"87",x"ee"),
  2115 => (x"f0",x"49",x"6a",x"4a"),
  2116 => (x"c6",x"f1",x"87",x"f0"),
  2117 => (x"c1",x"85",x"cb",x"87"),
  2118 => (x"ab",x"b7",x"c8",x"83"),
  2119 => (x"87",x"c7",x"ff",x"04"),
  2120 => (x"26",x"4d",x"26",x"26"),
  2121 => (x"26",x"4b",x"26",x"4c"),
  2122 => (x"4a",x"71",x"1e",x"4f"),
  2123 => (x"5a",x"ed",x"ec",x"c2"),
  2124 => (x"48",x"ed",x"ec",x"c2"),
  2125 => (x"fe",x"49",x"78",x"c7"),
  2126 => (x"4f",x"26",x"87",x"dd"),
  2127 => (x"71",x"1e",x"73",x"1e"),
  2128 => (x"aa",x"b7",x"c0",x"4a"),
  2129 => (x"c2",x"87",x"d3",x"03"),
  2130 => (x"05",x"bf",x"f8",x"d2"),
  2131 => (x"4b",x"c1",x"87",x"c4"),
  2132 => (x"4b",x"c0",x"87",x"c2"),
  2133 => (x"5b",x"fc",x"d2",x"c2"),
  2134 => (x"d2",x"c2",x"87",x"c4"),
  2135 => (x"d2",x"c2",x"5a",x"fc"),
  2136 => (x"c1",x"4a",x"bf",x"f8"),
  2137 => (x"a2",x"c0",x"c1",x"9a"),
  2138 => (x"87",x"e8",x"ec",x"49"),
  2139 => (x"d2",x"c2",x"48",x"fc"),
  2140 => (x"fe",x"78",x"bf",x"f8"),
  2141 => (x"71",x"1e",x"87",x"ef"),
  2142 => (x"1e",x"66",x"c4",x"4a"),
  2143 => (x"f9",x"ea",x"49",x"72"),
  2144 => (x"4f",x"26",x"26",x"87"),
  2145 => (x"48",x"d4",x"ff",x"1e"),
  2146 => (x"ff",x"78",x"ff",x"c3"),
  2147 => (x"e1",x"c0",x"48",x"d0"),
  2148 => (x"48",x"d4",x"ff",x"78"),
  2149 => (x"48",x"71",x"78",x"c1"),
  2150 => (x"d4",x"ff",x"30",x"c4"),
  2151 => (x"d0",x"ff",x"78",x"08"),
  2152 => (x"78",x"e0",x"c0",x"48"),
  2153 => (x"c2",x"1e",x"4f",x"26"),
  2154 => (x"49",x"bf",x"f8",x"d2"),
  2155 => (x"c2",x"87",x"f9",x"e6"),
  2156 => (x"e8",x"48",x"e1",x"ec"),
  2157 => (x"ec",x"c2",x"78",x"bf"),
  2158 => (x"bf",x"ec",x"48",x"dd"),
  2159 => (x"e1",x"ec",x"c2",x"78"),
  2160 => (x"c3",x"49",x"4a",x"bf"),
  2161 => (x"b7",x"c8",x"99",x"ff"),
  2162 => (x"71",x"48",x"72",x"2a"),
  2163 => (x"e9",x"ec",x"c2",x"b0"),
  2164 => (x"0e",x"4f",x"26",x"58"),
  2165 => (x"5d",x"5c",x"5b",x"5e"),
  2166 => (x"ff",x"4b",x"71",x"0e"),
  2167 => (x"ec",x"c2",x"87",x"c8"),
  2168 => (x"50",x"c0",x"48",x"dc"),
  2169 => (x"df",x"e6",x"49",x"73"),
  2170 => (x"4c",x"49",x"70",x"87"),
  2171 => (x"ee",x"cb",x"9c",x"c2"),
  2172 => (x"87",x"cc",x"cb",x"49"),
  2173 => (x"ec",x"c2",x"4d",x"70"),
  2174 => (x"05",x"bf",x"97",x"dc"),
  2175 => (x"d0",x"87",x"e2",x"c1"),
  2176 => (x"ec",x"c2",x"49",x"66"),
  2177 => (x"05",x"99",x"bf",x"e5"),
  2178 => (x"66",x"d4",x"87",x"d6"),
  2179 => (x"dd",x"ec",x"c2",x"49"),
  2180 => (x"cb",x"05",x"99",x"bf"),
  2181 => (x"e5",x"49",x"73",x"87"),
  2182 => (x"98",x"70",x"87",x"ee"),
  2183 => (x"87",x"c1",x"c1",x"02"),
  2184 => (x"c1",x"fe",x"4c",x"c1"),
  2185 => (x"ca",x"49",x"75",x"87"),
  2186 => (x"98",x"70",x"87",x"e2"),
  2187 => (x"c2",x"87",x"c6",x"02"),
  2188 => (x"c1",x"48",x"dc",x"ec"),
  2189 => (x"dc",x"ec",x"c2",x"50"),
  2190 => (x"c0",x"05",x"bf",x"97"),
  2191 => (x"ec",x"c2",x"87",x"e3"),
  2192 => (x"d0",x"49",x"bf",x"e5"),
  2193 => (x"ff",x"05",x"99",x"66"),
  2194 => (x"ec",x"c2",x"87",x"d6"),
  2195 => (x"d4",x"49",x"bf",x"dd"),
  2196 => (x"ff",x"05",x"99",x"66"),
  2197 => (x"49",x"73",x"87",x"ca"),
  2198 => (x"70",x"87",x"ed",x"e4"),
  2199 => (x"ff",x"fe",x"05",x"98"),
  2200 => (x"fa",x"48",x"74",x"87"),
  2201 => (x"5e",x"0e",x"87",x"fb"),
  2202 => (x"0e",x"5d",x"5c",x"5b"),
  2203 => (x"4d",x"c0",x"86",x"f8"),
  2204 => (x"7e",x"bf",x"ec",x"4c"),
  2205 => (x"c2",x"48",x"a6",x"c4"),
  2206 => (x"78",x"bf",x"e9",x"ec"),
  2207 => (x"1e",x"c0",x"1e",x"c1"),
  2208 => (x"ce",x"fd",x"49",x"c7"),
  2209 => (x"70",x"86",x"c8",x"87"),
  2210 => (x"87",x"cd",x"02",x"98"),
  2211 => (x"eb",x"fa",x"49",x"ff"),
  2212 => (x"49",x"da",x"c1",x"87"),
  2213 => (x"c1",x"87",x"f1",x"e3"),
  2214 => (x"dc",x"ec",x"c2",x"4d"),
  2215 => (x"cf",x"02",x"bf",x"97"),
  2216 => (x"f0",x"d2",x"c2",x"87"),
  2217 => (x"b9",x"c1",x"49",x"bf"),
  2218 => (x"59",x"f4",x"d2",x"c2"),
  2219 => (x"87",x"d4",x"fb",x"71"),
  2220 => (x"bf",x"e1",x"ec",x"c2"),
  2221 => (x"f8",x"d2",x"c2",x"4b"),
  2222 => (x"e9",x"c0",x"05",x"bf"),
  2223 => (x"49",x"fd",x"c3",x"87"),
  2224 => (x"c3",x"87",x"c5",x"e3"),
  2225 => (x"ff",x"e2",x"49",x"fa"),
  2226 => (x"c3",x"49",x"73",x"87"),
  2227 => (x"1e",x"71",x"99",x"ff"),
  2228 => (x"e1",x"fa",x"49",x"c0"),
  2229 => (x"c8",x"49",x"73",x"87"),
  2230 => (x"1e",x"71",x"29",x"b7"),
  2231 => (x"d5",x"fa",x"49",x"c1"),
  2232 => (x"c5",x"86",x"c8",x"87"),
  2233 => (x"ec",x"c2",x"87",x"f4"),
  2234 => (x"9b",x"4b",x"bf",x"e5"),
  2235 => (x"c2",x"87",x"dd",x"02"),
  2236 => (x"49",x"bf",x"f4",x"d2"),
  2237 => (x"70",x"87",x"d5",x"c7"),
  2238 => (x"87",x"c4",x"05",x"98"),
  2239 => (x"87",x"d2",x"4b",x"c0"),
  2240 => (x"c6",x"49",x"e0",x"c2"),
  2241 => (x"d2",x"c2",x"87",x"fa"),
  2242 => (x"87",x"c6",x"58",x"f8"),
  2243 => (x"48",x"f4",x"d2",x"c2"),
  2244 => (x"49",x"73",x"78",x"c0"),
  2245 => (x"cd",x"05",x"99",x"c2"),
  2246 => (x"49",x"eb",x"c3",x"87"),
  2247 => (x"70",x"87",x"e9",x"e1"),
  2248 => (x"02",x"99",x"c2",x"49"),
  2249 => (x"4c",x"fb",x"87",x"c2"),
  2250 => (x"99",x"c1",x"49",x"73"),
  2251 => (x"c3",x"87",x"cd",x"05"),
  2252 => (x"d3",x"e1",x"49",x"f4"),
  2253 => (x"c2",x"49",x"70",x"87"),
  2254 => (x"87",x"c2",x"02",x"99"),
  2255 => (x"49",x"73",x"4c",x"fa"),
  2256 => (x"cd",x"05",x"99",x"c8"),
  2257 => (x"49",x"f5",x"c3",x"87"),
  2258 => (x"70",x"87",x"fd",x"e0"),
  2259 => (x"02",x"99",x"c2",x"49"),
  2260 => (x"ec",x"c2",x"87",x"d5"),
  2261 => (x"ca",x"02",x"bf",x"ed"),
  2262 => (x"88",x"c1",x"48",x"87"),
  2263 => (x"58",x"f1",x"ec",x"c2"),
  2264 => (x"ff",x"87",x"c2",x"c0"),
  2265 => (x"73",x"4d",x"c1",x"4c"),
  2266 => (x"05",x"99",x"c4",x"49"),
  2267 => (x"f2",x"c3",x"87",x"cd"),
  2268 => (x"87",x"d4",x"e0",x"49"),
  2269 => (x"99",x"c2",x"49",x"70"),
  2270 => (x"c2",x"87",x"dc",x"02"),
  2271 => (x"7e",x"bf",x"ed",x"ec"),
  2272 => (x"a8",x"b7",x"c7",x"48"),
  2273 => (x"87",x"cb",x"c0",x"03"),
  2274 => (x"80",x"c1",x"48",x"6e"),
  2275 => (x"58",x"f1",x"ec",x"c2"),
  2276 => (x"fe",x"87",x"c2",x"c0"),
  2277 => (x"c3",x"4d",x"c1",x"4c"),
  2278 => (x"df",x"ff",x"49",x"fd"),
  2279 => (x"49",x"70",x"87",x"ea"),
  2280 => (x"d5",x"02",x"99",x"c2"),
  2281 => (x"ed",x"ec",x"c2",x"87"),
  2282 => (x"c9",x"c0",x"02",x"bf"),
  2283 => (x"ed",x"ec",x"c2",x"87"),
  2284 => (x"c0",x"78",x"c0",x"48"),
  2285 => (x"4c",x"fd",x"87",x"c2"),
  2286 => (x"fa",x"c3",x"4d",x"c1"),
  2287 => (x"c7",x"df",x"ff",x"49"),
  2288 => (x"c2",x"49",x"70",x"87"),
  2289 => (x"d9",x"c0",x"02",x"99"),
  2290 => (x"ed",x"ec",x"c2",x"87"),
  2291 => (x"b7",x"c7",x"48",x"bf"),
  2292 => (x"c9",x"c0",x"03",x"a8"),
  2293 => (x"ed",x"ec",x"c2",x"87"),
  2294 => (x"c0",x"78",x"c7",x"48"),
  2295 => (x"4c",x"fc",x"87",x"c2"),
  2296 => (x"b7",x"c0",x"4d",x"c1"),
  2297 => (x"d3",x"c0",x"03",x"ac"),
  2298 => (x"48",x"66",x"c4",x"87"),
  2299 => (x"70",x"80",x"d8",x"c1"),
  2300 => (x"02",x"bf",x"6e",x"7e"),
  2301 => (x"4b",x"87",x"c5",x"c0"),
  2302 => (x"0f",x"73",x"49",x"74"),
  2303 => (x"f0",x"c3",x"1e",x"c0"),
  2304 => (x"49",x"da",x"c1",x"1e"),
  2305 => (x"c8",x"87",x"cc",x"f7"),
  2306 => (x"02",x"98",x"70",x"86"),
  2307 => (x"c2",x"87",x"d8",x"c0"),
  2308 => (x"7e",x"bf",x"ed",x"ec"),
  2309 => (x"91",x"cb",x"49",x"6e"),
  2310 => (x"71",x"4a",x"66",x"c4"),
  2311 => (x"c0",x"02",x"6a",x"82"),
  2312 => (x"6e",x"4b",x"87",x"c5"),
  2313 => (x"75",x"0f",x"73",x"49"),
  2314 => (x"c8",x"c0",x"02",x"9d"),
  2315 => (x"ed",x"ec",x"c2",x"87"),
  2316 => (x"e2",x"f2",x"49",x"bf"),
  2317 => (x"fc",x"d2",x"c2",x"87"),
  2318 => (x"dd",x"c0",x"02",x"bf"),
  2319 => (x"cb",x"c2",x"49",x"87"),
  2320 => (x"02",x"98",x"70",x"87"),
  2321 => (x"c2",x"87",x"d3",x"c0"),
  2322 => (x"49",x"bf",x"ed",x"ec"),
  2323 => (x"c0",x"87",x"c8",x"f2"),
  2324 => (x"87",x"e8",x"f3",x"49"),
  2325 => (x"48",x"fc",x"d2",x"c2"),
  2326 => (x"8e",x"f8",x"78",x"c0"),
  2327 => (x"0e",x"87",x"c2",x"f3"),
  2328 => (x"5d",x"5c",x"5b",x"5e"),
  2329 => (x"4c",x"71",x"1e",x"0e"),
  2330 => (x"bf",x"e9",x"ec",x"c2"),
  2331 => (x"a1",x"cd",x"c1",x"49"),
  2332 => (x"81",x"d1",x"c1",x"4d"),
  2333 => (x"9c",x"74",x"7e",x"69"),
  2334 => (x"c4",x"87",x"cf",x"02"),
  2335 => (x"7b",x"74",x"4b",x"a5"),
  2336 => (x"bf",x"e9",x"ec",x"c2"),
  2337 => (x"87",x"e1",x"f2",x"49"),
  2338 => (x"9c",x"74",x"7b",x"6e"),
  2339 => (x"c0",x"87",x"c4",x"05"),
  2340 => (x"c1",x"87",x"c2",x"4b"),
  2341 => (x"f2",x"49",x"73",x"4b"),
  2342 => (x"66",x"d4",x"87",x"e2"),
  2343 => (x"49",x"87",x"c7",x"02"),
  2344 => (x"4a",x"70",x"87",x"de"),
  2345 => (x"4a",x"c0",x"87",x"c2"),
  2346 => (x"5a",x"c0",x"d3",x"c2"),
  2347 => (x"87",x"f1",x"f1",x"26"),
  2348 => (x"00",x"00",x"00",x"00"),
  2349 => (x"00",x"00",x"00",x"00"),
  2350 => (x"00",x"00",x"00",x"00"),
  2351 => (x"00",x"00",x"00",x"00"),
  2352 => (x"ff",x"4a",x"71",x"1e"),
  2353 => (x"72",x"49",x"bf",x"c8"),
  2354 => (x"4f",x"26",x"48",x"a1"),
  2355 => (x"bf",x"c8",x"ff",x"1e"),
  2356 => (x"c0",x"c0",x"fe",x"89"),
  2357 => (x"a9",x"c0",x"c0",x"c0"),
  2358 => (x"c0",x"87",x"c4",x"01"),
  2359 => (x"c1",x"87",x"c2",x"4a"),
  2360 => (x"26",x"48",x"72",x"4a"),
  2361 => (x"5b",x"5e",x"0e",x"4f"),
  2362 => (x"71",x"0e",x"5d",x"5c"),
  2363 => (x"4c",x"d4",x"ff",x"4b"),
  2364 => (x"c0",x"48",x"66",x"d0"),
  2365 => (x"ff",x"49",x"d6",x"78"),
  2366 => (x"c3",x"87",x"c5",x"dc"),
  2367 => (x"49",x"6c",x"7c",x"ff"),
  2368 => (x"71",x"99",x"ff",x"c3"),
  2369 => (x"f0",x"c3",x"49",x"4d"),
  2370 => (x"a9",x"e0",x"c1",x"99"),
  2371 => (x"c3",x"87",x"cb",x"05"),
  2372 => (x"48",x"6c",x"7c",x"ff"),
  2373 => (x"66",x"d0",x"98",x"c3"),
  2374 => (x"ff",x"c3",x"78",x"08"),
  2375 => (x"49",x"4a",x"6c",x"7c"),
  2376 => (x"ff",x"c3",x"31",x"c8"),
  2377 => (x"71",x"4a",x"6c",x"7c"),
  2378 => (x"c8",x"49",x"72",x"b2"),
  2379 => (x"7c",x"ff",x"c3",x"31"),
  2380 => (x"b2",x"71",x"4a",x"6c"),
  2381 => (x"31",x"c8",x"49",x"72"),
  2382 => (x"6c",x"7c",x"ff",x"c3"),
  2383 => (x"ff",x"b2",x"71",x"4a"),
  2384 => (x"e0",x"c0",x"48",x"d0"),
  2385 => (x"02",x"9b",x"73",x"78"),
  2386 => (x"7b",x"72",x"87",x"c2"),
  2387 => (x"4d",x"26",x"48",x"75"),
  2388 => (x"4b",x"26",x"4c",x"26"),
  2389 => (x"26",x"1e",x"4f",x"26"),
  2390 => (x"5b",x"5e",x"0e",x"4f"),
  2391 => (x"86",x"f8",x"0e",x"5c"),
  2392 => (x"a6",x"c8",x"1e",x"76"),
  2393 => (x"87",x"fd",x"fd",x"49"),
  2394 => (x"4b",x"70",x"86",x"c4"),
  2395 => (x"a8",x"c4",x"48",x"6e"),
  2396 => (x"87",x"f0",x"c2",x"03"),
  2397 => (x"f0",x"c3",x"4a",x"73"),
  2398 => (x"aa",x"d0",x"c1",x"9a"),
  2399 => (x"c1",x"87",x"c7",x"02"),
  2400 => (x"c2",x"05",x"aa",x"e0"),
  2401 => (x"49",x"73",x"87",x"de"),
  2402 => (x"c3",x"02",x"99",x"c8"),
  2403 => (x"87",x"c6",x"ff",x"87"),
  2404 => (x"9c",x"c3",x"4c",x"73"),
  2405 => (x"c1",x"05",x"ac",x"c2"),
  2406 => (x"66",x"c4",x"87",x"c2"),
  2407 => (x"71",x"31",x"c9",x"49"),
  2408 => (x"4a",x"66",x"c4",x"1e"),
  2409 => (x"ec",x"c2",x"92",x"d4"),
  2410 => (x"81",x"72",x"49",x"f1"),
  2411 => (x"87",x"d9",x"d0",x"fe"),
  2412 => (x"d9",x"ff",x"49",x"d8"),
  2413 => (x"c0",x"c8",x"87",x"ca"),
  2414 => (x"ce",x"db",x"c2",x"1e"),
  2415 => (x"dd",x"ec",x"fd",x"49"),
  2416 => (x"48",x"d0",x"ff",x"87"),
  2417 => (x"c2",x"78",x"e0",x"c0"),
  2418 => (x"cc",x"1e",x"ce",x"db"),
  2419 => (x"92",x"d4",x"4a",x"66"),
  2420 => (x"49",x"f1",x"ec",x"c2"),
  2421 => (x"ce",x"fe",x"81",x"72"),
  2422 => (x"86",x"cc",x"87",x"e1"),
  2423 => (x"c1",x"05",x"ac",x"c1"),
  2424 => (x"66",x"c4",x"87",x"c2"),
  2425 => (x"71",x"31",x"c9",x"49"),
  2426 => (x"4a",x"66",x"c4",x"1e"),
  2427 => (x"ec",x"c2",x"92",x"d4"),
  2428 => (x"81",x"72",x"49",x"f1"),
  2429 => (x"87",x"d1",x"cf",x"fe"),
  2430 => (x"1e",x"ce",x"db",x"c2"),
  2431 => (x"d4",x"4a",x"66",x"c8"),
  2432 => (x"f1",x"ec",x"c2",x"92"),
  2433 => (x"fe",x"81",x"72",x"49"),
  2434 => (x"d7",x"87",x"e2",x"cc"),
  2435 => (x"ef",x"d7",x"ff",x"49"),
  2436 => (x"1e",x"c0",x"c8",x"87"),
  2437 => (x"49",x"ce",x"db",x"c2"),
  2438 => (x"87",x"db",x"ea",x"fd"),
  2439 => (x"d0",x"ff",x"86",x"cc"),
  2440 => (x"78",x"e0",x"c0",x"48"),
  2441 => (x"e7",x"fc",x"8e",x"f8"),
  2442 => (x"5b",x"5e",x"0e",x"87"),
  2443 => (x"71",x"0e",x"5d",x"5c"),
  2444 => (x"4c",x"d4",x"ff",x"4a"),
  2445 => (x"c3",x"4d",x"66",x"d0"),
  2446 => (x"c5",x"06",x"ad",x"b7"),
  2447 => (x"c1",x"48",x"c0",x"87"),
  2448 => (x"1e",x"72",x"87",x"e1"),
  2449 => (x"93",x"d4",x"4b",x"75"),
  2450 => (x"83",x"f1",x"ec",x"c2"),
  2451 => (x"c6",x"fe",x"49",x"73"),
  2452 => (x"83",x"c8",x"87",x"e7"),
  2453 => (x"d0",x"ff",x"4b",x"6b"),
  2454 => (x"78",x"e1",x"c8",x"48"),
  2455 => (x"48",x"73",x"7c",x"dd"),
  2456 => (x"70",x"98",x"ff",x"c3"),
  2457 => (x"c8",x"49",x"73",x"7c"),
  2458 => (x"48",x"71",x"29",x"b7"),
  2459 => (x"70",x"98",x"ff",x"c3"),
  2460 => (x"d0",x"49",x"73",x"7c"),
  2461 => (x"48",x"71",x"29",x"b7"),
  2462 => (x"70",x"98",x"ff",x"c3"),
  2463 => (x"d8",x"48",x"73",x"7c"),
  2464 => (x"7c",x"70",x"28",x"b7"),
  2465 => (x"7c",x"7c",x"7c",x"c0"),
  2466 => (x"7c",x"7c",x"7c",x"7c"),
  2467 => (x"7c",x"7c",x"7c",x"7c"),
  2468 => (x"48",x"d0",x"ff",x"7c"),
  2469 => (x"75",x"78",x"e0",x"c0"),
  2470 => (x"ff",x"49",x"dc",x"1e"),
  2471 => (x"c8",x"87",x"c6",x"d6"),
  2472 => (x"fa",x"48",x"73",x"86"),
  2473 => (x"fa",x"48",x"87",x"e8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

