library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4eec287",
    12 => x"86c0c84e",
    13 => x"49c4eec2",
    14 => x"48e8dac2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e9e2",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfe8da",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dac21e73",
   183 => x"78c148e8",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"ecdac287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58f0dac2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49f0dac2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97f0da",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97f7da",
   291 => x"c231d049",
   292 => x"bf97f8da",
   293 => x"7232c84a",
   294 => x"f9dac2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dac287e7",
   300 => x"49bf97f9",
   301 => x"99c631c1",
   302 => x"97fadac2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97f5da",
   306 => x"9dcf4d4a",
   307 => x"97f6dac2",
   308 => x"9ac34abf",
   309 => x"dac232ca",
   310 => x"4bbf97f7",
   311 => x"b27333c2",
   312 => x"97f8dac2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e3c286f8",
   329 => x"78c048d6",
   330 => x"1ecedbc2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"e2f2c07e",
   337 => x"dcc249bf",
   338 => x"c8714ac4",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfdef2",
   343 => x"4ae0dcc2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e2c287fd",
   349 => x"c24dbfd4",
   350 => x"bf9fcce3",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"d4e2c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"dbc287e3",
   359 => x"49751ece",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfdef2",
   365 => x"4ae0dcc2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148d6e3",
   370 => x"c087da78",
   371 => x"49bfe2f2",
   372 => x"4ac4dcc2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"cce3c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e3c287cd",
   381 => x"49bf97cd",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97cedbc2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97d9dbc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97dadb",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97dbdbc2",
   400 => x"e3c248bf",
   401 => x"4c7058d2",
   402 => x"c288c148",
   403 => x"c258d6e3",
   404 => x"bf97dcdb",
   405 => x"c2817549",
   406 => x"bf97dddb",
   407 => x"7232c84a",
   408 => x"e7c27ea1",
   409 => x"786e48e3",
   410 => x"97dedbc2",
   411 => x"a6c848bf",
   412 => x"d6e3c258",
   413 => x"cfc202bf",
   414 => x"def2c087",
   415 => x"dcc249bf",
   416 => x"c8714ae0",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbfcee3",
   422 => x"5cf7e7c2",
   423 => x"97f3dbc2",
   424 => x"31c849bf",
   425 => x"97f2dbc2",
   426 => x"49a14abf",
   427 => x"97f4dbc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97f5db",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"e3e7c291",
   434 => x"e7c281bf",
   435 => x"dbc259eb",
   436 => x"4abf97fb",
   437 => x"dbc232c8",
   438 => x"4bbf97fa",
   439 => x"dbc24aa2",
   440 => x"4bbf97fc",
   441 => x"a27333d0",
   442 => x"fddbc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e7c24aa2",
   446 => x"8ac25aef",
   447 => x"e7c29274",
   448 => x"a17248ef",
   449 => x"87c1c178",
   450 => x"97e0dbc2",
   451 => x"31c849bf",
   452 => x"97dfdbc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259f7e7",
   457 => x"bf97e5db",
   458 => x"c232c84a",
   459 => x"bf97e4db",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5af3e7c2",
   463 => x"48ebe7c2",
   464 => x"e7c278c0",
   465 => x"a17248e7",
   466 => x"f7e7c278",
   467 => x"ebe7c248",
   468 => x"e7c278bf",
   469 => x"e7c248fb",
   470 => x"c278bfef",
   471 => x"02bfd6e3",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bff3e7c2",
   476 => x"7030c448",
   477 => x"dae3c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfd6e3",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e7c29dff",
   491 => x"c083bfe3",
   492 => x"abbfdaf2",
   493 => x"c087d902",
   494 => x"c25bdef2",
   495 => x"731ecedb",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfd6e3c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981cedb",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"cedbc291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c1c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087eac2",
   521 => x"4949c11e",
   522 => x"c487d6ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4adee3c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d4c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cfc102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfd6e3",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"496e7ec0",
   556 => x"bf66c448",
   557 => x"0866c480",
   558 => x"cc7cc078",
   559 => x"66c449a4",
   560 => x"a4d079bf",
   561 => x"c179c049",
   562 => x"c087c248",
   563 => x"fa8ef848",
   564 => x"5e0e87ed",
   565 => x"0e5d5c5b",
   566 => x"029c4c71",
   567 => x"c887cbc1",
   568 => x"026949a4",
   569 => x"d087c3c1",
   570 => x"496c4a66",
   571 => x"7248a6d0",
   572 => x"b94d78a1",
   573 => x"bfd2e3c2",
   574 => x"72baff4a",
   575 => x"02997199",
   576 => x"c487e4c0",
   577 => x"496b4ba4",
   578 => x"7087fcf9",
   579 => x"cee3c27b",
   580 => x"816c49bf",
   581 => x"b9757c71",
   582 => x"bfd2e3c2",
   583 => x"72baff4a",
   584 => x"05997199",
   585 => x"d087dcff",
   586 => x"d2f97c66",
   587 => x"1e731e87",
   588 => x"029b4b71",
   589 => x"a3c887c7",
   590 => x"c5056949",
   591 => x"c048c087",
   592 => x"e7c287f6",
   593 => x"c449bfe7",
   594 => x"4a6a4aa3",
   595 => x"e3c28ac2",
   596 => x"7292bfce",
   597 => x"e3c249a1",
   598 => x"6b4abfd2",
   599 => x"49a1729a",
   600 => x"59def2c0",
   601 => x"711e66c8",
   602 => x"c487e4ea",
   603 => x"05987086",
   604 => x"48c087c4",
   605 => x"48c187c2",
   606 => x"1e87c8f8",
   607 => x"4b711e73",
   608 => x"87c7029b",
   609 => x"6949a3c8",
   610 => x"c087c505",
   611 => x"87f6c048",
   612 => x"bfe7e7c2",
   613 => x"4aa3c449",
   614 => x"8ac24a6a",
   615 => x"bfcee3c2",
   616 => x"49a17292",
   617 => x"bfd2e3c2",
   618 => x"729a6b4a",
   619 => x"f2c049a1",
   620 => x"66c859de",
   621 => x"cfe6711e",
   622 => x"7086c487",
   623 => x"87c40598",
   624 => x"87c248c0",
   625 => x"faf648c1",
   626 => x"5b5e0e87",
   627 => x"1e0e5d5c",
   628 => x"66d44b71",
   629 => x"029b734d",
   630 => x"c887ccc1",
   631 => x"026949a3",
   632 => x"d087c4c1",
   633 => x"e3c24ca3",
   634 => x"ff49bfd2",
   635 => x"994a6cb9",
   636 => x"a966d47e",
   637 => x"c087cd06",
   638 => x"a3cc7c7b",
   639 => x"49a3c44a",
   640 => x"87ca796a",
   641 => x"c0f84972",
   642 => x"4d66d499",
   643 => x"49758d71",
   644 => x"1e7129c9",
   645 => x"f9fa4973",
   646 => x"cedbc287",
   647 => x"fc49731e",
   648 => x"86c887cb",
   649 => x"267c66d4",
   650 => x"1e87d4f5",
   651 => x"4b711e73",
   652 => x"e4c0029b",
   653 => x"fbe7c287",
   654 => x"c24a735b",
   655 => x"cee3c28a",
   656 => x"c29249bf",
   657 => x"48bfe7e7",
   658 => x"e7c28072",
   659 => x"487158ff",
   660 => x"e3c230c4",
   661 => x"edc058de",
   662 => x"f7e7c287",
   663 => x"ebe7c248",
   664 => x"e7c278bf",
   665 => x"e7c248fb",
   666 => x"c278bfef",
   667 => x"02bfd6e3",
   668 => x"e3c287c9",
   669 => x"c449bfce",
   670 => x"c287c731",
   671 => x"49bff3e7",
   672 => x"e3c231c4",
   673 => x"faf359de",
   674 => x"5b5e0e87",
   675 => x"4a710e5c",
   676 => x"9a724bc0",
   677 => x"87e1c002",
   678 => x"9f49a2da",
   679 => x"e3c24b69",
   680 => x"cf02bfd6",
   681 => x"49a2d487",
   682 => x"4c49699f",
   683 => x"9cffffc0",
   684 => x"87c234d0",
   685 => x"49744cc0",
   686 => x"fd4973b3",
   687 => x"c0f387ed",
   688 => x"5b5e0e87",
   689 => x"f40e5d5c",
   690 => x"c04a7186",
   691 => x"029a727e",
   692 => x"dbc287d8",
   693 => x"78c048ca",
   694 => x"48c2dbc2",
   695 => x"bffbe7c2",
   696 => x"c6dbc278",
   697 => x"f7e7c248",
   698 => x"e3c278bf",
   699 => x"50c048eb",
   700 => x"bfdae3c2",
   701 => x"cadbc249",
   702 => x"aa714abf",
   703 => x"87c9c403",
   704 => x"99cf4972",
   705 => x"87e9c005",
   706 => x"48daf2c0",
   707 => x"bfc2dbc2",
   708 => x"cedbc278",
   709 => x"c2dbc21e",
   710 => x"dbc249bf",
   711 => x"a1c148c2",
   712 => x"eae37178",
   713 => x"c086c487",
   714 => x"c248d6f2",
   715 => x"cc78cedb",
   716 => x"d6f2c087",
   717 => x"e0c048bf",
   718 => x"daf2c080",
   719 => x"cadbc258",
   720 => x"80c148bf",
   721 => x"58cedbc2",
   722 => x"000c9627",
   723 => x"bf97bf00",
   724 => x"c2029d4d",
   725 => x"e5c387e3",
   726 => x"dcc202ad",
   727 => x"d6f2c087",
   728 => x"a3cb4bbf",
   729 => x"cf4c1149",
   730 => x"d2c105ac",
   731 => x"df497587",
   732 => x"cd89c199",
   733 => x"dee3c291",
   734 => x"4aa3c181",
   735 => x"a3c35112",
   736 => x"c551124a",
   737 => x"51124aa3",
   738 => x"124aa3c7",
   739 => x"4aa3c951",
   740 => x"a3ce5112",
   741 => x"d051124a",
   742 => x"51124aa3",
   743 => x"124aa3d2",
   744 => x"4aa3d451",
   745 => x"a3d65112",
   746 => x"d851124a",
   747 => x"51124aa3",
   748 => x"124aa3dc",
   749 => x"4aa3de51",
   750 => x"7ec15112",
   751 => x"7487fac0",
   752 => x"0599c849",
   753 => x"7487ebc0",
   754 => x"0599d049",
   755 => x"66dc87d1",
   756 => x"87cbc002",
   757 => x"66dc4973",
   758 => x"0298700f",
   759 => x"6e87d3c0",
   760 => x"87c6c005",
   761 => x"48dee3c2",
   762 => x"f2c050c0",
   763 => x"c248bfd6",
   764 => x"e3c287df",
   765 => x"50c048eb",
   766 => x"dae3c27e",
   767 => x"dbc249bf",
   768 => x"714abfca",
   769 => x"f7fb04aa",
   770 => x"fbe7c287",
   771 => x"c8c005bf",
   772 => x"d6e3c287",
   773 => x"f6c102bf",
   774 => x"c6dbc287",
   775 => x"e6ed49bf",
   776 => x"cadbc287",
   777 => x"48a6c458",
   778 => x"bfc6dbc2",
   779 => x"d6e3c278",
   780 => x"d8c002bf",
   781 => x"4966c487",
   782 => x"ffffffcf",
   783 => x"02a999f8",
   784 => x"c087c5c0",
   785 => x"87e1c04c",
   786 => x"dcc04cc1",
   787 => x"4966c487",
   788 => x"99f8ffcf",
   789 => x"c8c002a9",
   790 => x"48a6c887",
   791 => x"c5c078c0",
   792 => x"48a6c887",
   793 => x"66c878c1",
   794 => x"059c744c",
   795 => x"c487e0c0",
   796 => x"89c24966",
   797 => x"bfcee3c2",
   798 => x"e7c2914a",
   799 => x"c24abfe7",
   800 => x"7248c2db",
   801 => x"dbc278a1",
   802 => x"78c048ca",
   803 => x"c087e1f9",
   804 => x"eb8ef448",
   805 => x"000087e9",
   806 => x"ffff0000",
   807 => x"0ca6ffff",
   808 => x"0caf0000",
   809 => x"41460000",
   810 => x"20323354",
   811 => x"46002020",
   812 => x"36315441",
   813 => x"00202020",
   814 => x"48d4ff1e",
   815 => x"6878ffc3",
   816 => x"1e4f2648",
   817 => x"c348d4ff",
   818 => x"d0ff78ff",
   819 => x"78e1c048",
   820 => x"d448d4ff",
   821 => x"ffe7c278",
   822 => x"bfd4ff48",
   823 => x"1e4f2650",
   824 => x"c048d0ff",
   825 => x"4f2678e0",
   826 => x"87ccff1e",
   827 => x"02994970",
   828 => x"fbc087c6",
   829 => x"87f105a9",
   830 => x"4f264871",
   831 => x"5c5b5e0e",
   832 => x"c04b710e",
   833 => x"87f0fe4c",
   834 => x"02994970",
   835 => x"c087f9c0",
   836 => x"c002a9ec",
   837 => x"fbc087f2",
   838 => x"ebc002a9",
   839 => x"b766cc87",
   840 => x"87c703ac",
   841 => x"c20266d0",
   842 => x"71537187",
   843 => x"87c20299",
   844 => x"c3fe84c1",
   845 => x"99497087",
   846 => x"c087cd02",
   847 => x"c702a9ec",
   848 => x"a9fbc087",
   849 => x"87d5ff05",
   850 => x"c30266d0",
   851 => x"7b97c087",
   852 => x"05a9ecc0",
   853 => x"4a7487c4",
   854 => x"4a7487c5",
   855 => x"728a0ac0",
   856 => x"2687c248",
   857 => x"264c264d",
   858 => x"1e4f264b",
   859 => x"7087c9fd",
   860 => x"aaf0c04a",
   861 => x"c087c904",
   862 => x"c301aaf9",
   863 => x"8af0c087",
   864 => x"04aac1c1",
   865 => x"dac187c9",
   866 => x"87c301aa",
   867 => x"728af7c0",
   868 => x"0e4f2648",
   869 => x"5d5c5b5e",
   870 => x"7186f80e",
   871 => x"fc7ec04c",
   872 => x"4bc087e1",
   873 => x"97c0f9c0",
   874 => x"a9c049bf",
   875 => x"fc87cf04",
   876 => x"83c187f6",
   877 => x"97c0f9c0",
   878 => x"06ab49bf",
   879 => x"f9c087f1",
   880 => x"02bf97c0",
   881 => x"effb87cf",
   882 => x"99497087",
   883 => x"c087c602",
   884 => x"f105a9ec",
   885 => x"fb4bc087",
   886 => x"4d7087de",
   887 => x"c887d9fb",
   888 => x"d3fb58a6",
   889 => x"c14a7087",
   890 => x"49a4c883",
   891 => x"ad496997",
   892 => x"c087c702",
   893 => x"c005adff",
   894 => x"a4c987e7",
   895 => x"49699749",
   896 => x"02a966c4",
   897 => x"c04887c7",
   898 => x"d405a8ff",
   899 => x"49a4ca87",
   900 => x"aa496997",
   901 => x"c087c602",
   902 => x"c405aaff",
   903 => x"d07ec187",
   904 => x"adecc087",
   905 => x"c087c602",
   906 => x"c405adfb",
   907 => x"c14bc087",
   908 => x"fe026e7e",
   909 => x"e6fa87e1",
   910 => x"f8487387",
   911 => x"87e3fc8e",
   912 => x"5b5e0e00",
   913 => x"f40e5d5c",
   914 => x"ff7e7186",
   915 => x"1e6e4bd4",
   916 => x"49c4e8c2",
   917 => x"c487e2e6",
   918 => x"02987086",
   919 => x"c487f5c4",
   920 => x"e4c148a6",
   921 => x"6e78bfcc",
   922 => x"87e7fc49",
   923 => x"7058a6cc",
   924 => x"87c50598",
   925 => x"c148a6c8",
   926 => x"48d0ff78",
   927 => x"d5c178c5",
   928 => x"4966c87b",
   929 => x"31c689c1",
   930 => x"97cae4c1",
   931 => x"71484abf",
   932 => x"ff7b70b0",
   933 => x"78c448d0",
   934 => x"d6c178c5",
   935 => x"6e4dc07b",
   936 => x"11817549",
   937 => x"cb85c17b",
   938 => x"f204adb7",
   939 => x"c34dcc87",
   940 => x"85c17bff",
   941 => x"adb7e0c0",
   942 => x"ff87f404",
   943 => x"78c448d0",
   944 => x"c57bffc3",
   945 => x"7bd3c178",
   946 => x"78c47bc1",
   947 => x"b7c04866",
   948 => x"eec206a8",
   949 => x"cce8c287",
   950 => x"66c44cbf",
   951 => x"c8887448",
   952 => x"9c7458a6",
   953 => x"87f7c102",
   954 => x"7ecedbc2",
   955 => x"8c4dc0c8",
   956 => x"03acb7c0",
   957 => x"c0c887c6",
   958 => x"4cc04da4",
   959 => x"97ffe7c2",
   960 => x"99d049bf",
   961 => x"c087d002",
   962 => x"c4e8c21e",
   963 => x"87dde849",
   964 => x"4a7086c4",
   965 => x"c287edc0",
   966 => x"c21ecedb",
   967 => x"e849c4e8",
   968 => x"86c487cb",
   969 => x"d0ff4a70",
   970 => x"78c5c848",
   971 => x"6e7bd4c1",
   972 => x"6e7bbf97",
   973 => x"7080c148",
   974 => x"058dc17e",
   975 => x"ff87f0ff",
   976 => x"78c448d0",
   977 => x"c5059a72",
   978 => x"c148c087",
   979 => x"1ec187c8",
   980 => x"49c4e8c2",
   981 => x"c487fbe5",
   982 => x"059c7486",
   983 => x"c487c9fe",
   984 => x"b7c04866",
   985 => x"87d106a8",
   986 => x"48c4e8c2",
   987 => x"80d078c0",
   988 => x"80f478c0",
   989 => x"bfd0e8c2",
   990 => x"4866c478",
   991 => x"01a8b7c0",
   992 => x"ff87d2fd",
   993 => x"78c548d0",
   994 => x"c07bd3c1",
   995 => x"c178c47b",
   996 => x"87c2c048",
   997 => x"8ef448c0",
   998 => x"4c264d26",
   999 => x"4f264b26",
  1000 => x"5c5b5e0e",
  1001 => x"711e0e5d",
  1002 => x"4d4cc04b",
  1003 => x"e8c004ab",
  1004 => x"d3f6c087",
  1005 => x"029d751e",
  1006 => x"4ac087c4",
  1007 => x"4ac187c2",
  1008 => x"fceb4972",
  1009 => x"7086c487",
  1010 => x"6e84c17e",
  1011 => x"7387c205",
  1012 => x"7385c14c",
  1013 => x"d8ff06ac",
  1014 => x"26486e87",
  1015 => x"0e87f9fe",
  1016 => x"0e5c5b5e",
  1017 => x"66cc4b71",
  1018 => x"4c87d802",
  1019 => x"028cf0c0",
  1020 => x"4a7487d8",
  1021 => x"d1028ac1",
  1022 => x"cd028a87",
  1023 => x"c9028a87",
  1024 => x"7387d987",
  1025 => x"87f9f849",
  1026 => x"1e7487d2",
  1027 => x"d8c149c0",
  1028 => x"1e7487d7",
  1029 => x"d8c14973",
  1030 => x"86c887cf",
  1031 => x"0e87fbfd",
  1032 => x"5d5c5b5e",
  1033 => x"4c711e0e",
  1034 => x"c291de49",
  1035 => x"714dece8",
  1036 => x"026d9785",
  1037 => x"c287dcc1",
  1038 => x"49bfd8e8",
  1039 => x"fd718174",
  1040 => x"7e7087de",
  1041 => x"c0029848",
  1042 => x"e8c287f2",
  1043 => x"4a704be0",
  1044 => x"c1ff49cb",
  1045 => x"4b7487d1",
  1046 => x"e4c193cb",
  1047 => x"83c483de",
  1048 => x"7bd7c2c1",
  1049 => x"c1c14974",
  1050 => x"7b7587ed",
  1051 => x"97cbe4c1",
  1052 => x"c21e49bf",
  1053 => x"fd49e0e8",
  1054 => x"86c487e5",
  1055 => x"c1c14974",
  1056 => x"49c087d5",
  1057 => x"87f4c2c1",
  1058 => x"48c0e8c2",
  1059 => x"49c178c0",
  1060 => x"2687fbdd",
  1061 => x"4c87c1fc",
  1062 => x"6964616f",
  1063 => x"2e2e676e",
  1064 => x"731e002e",
  1065 => x"494a711e",
  1066 => x"bfd8e8c2",
  1067 => x"effb7181",
  1068 => x"9b4b7087",
  1069 => x"4987c402",
  1070 => x"c287cee7",
  1071 => x"c048d8e8",
  1072 => x"dd49c178",
  1073 => x"d3fb87c8",
  1074 => x"49c01e87",
  1075 => x"87ecc1c1",
  1076 => x"711e4f26",
  1077 => x"91cb494a",
  1078 => x"81dee4c1",
  1079 => x"481181c8",
  1080 => x"58c4e8c2",
  1081 => x"48d8e8c2",
  1082 => x"49c178c0",
  1083 => x"2687dfdc",
  1084 => x"99711e4f",
  1085 => x"c187d202",
  1086 => x"c048f3e5",
  1087 => x"c180f750",
  1088 => x"c140d2c3",
  1089 => x"ce78d7e4",
  1090 => x"efe5c187",
  1091 => x"d0e4c148",
  1092 => x"c180fc78",
  1093 => x"2678c9c3",
  1094 => x"5b5e0e4f",
  1095 => x"f40e5d5c",
  1096 => x"cedbc286",
  1097 => x"c44cc04d",
  1098 => x"78c048a6",
  1099 => x"bfd8e8c2",
  1100 => x"06a8c048",
  1101 => x"c287c0c1",
  1102 => x"9848cedb",
  1103 => x"87f7c002",
  1104 => x"1ed3f6c0",
  1105 => x"c70266c8",
  1106 => x"48a6c487",
  1107 => x"87c578c0",
  1108 => x"c148a6c4",
  1109 => x"4966c478",
  1110 => x"c487e6e5",
  1111 => x"c14d7086",
  1112 => x"4866c484",
  1113 => x"a6c880c1",
  1114 => x"d8e8c258",
  1115 => x"c603acbf",
  1116 => x"059d7587",
  1117 => x"c087c9ff",
  1118 => x"029d754c",
  1119 => x"c087dcc3",
  1120 => x"c81ed3f6",
  1121 => x"87c70266",
  1122 => x"c048a6cc",
  1123 => x"cc87c578",
  1124 => x"78c148a6",
  1125 => x"e44966cc",
  1126 => x"86c487e7",
  1127 => x"98487e70",
  1128 => x"87e4c202",
  1129 => x"9781cb49",
  1130 => x"99d04969",
  1131 => x"87d4c102",
  1132 => x"91cb4974",
  1133 => x"81dee4c1",
  1134 => x"79e2c2c1",
  1135 => x"ffc381c8",
  1136 => x"de497451",
  1137 => x"ece8c291",
  1138 => x"c285714d",
  1139 => x"c17d97c1",
  1140 => x"e0c049a5",
  1141 => x"dee3c251",
  1142 => x"d202bf97",
  1143 => x"c284c187",
  1144 => x"e3c24ba5",
  1145 => x"49db4ade",
  1146 => x"87fbfafe",
  1147 => x"cd87d9c1",
  1148 => x"51c049a5",
  1149 => x"a5c284c1",
  1150 => x"cb4a6e4b",
  1151 => x"e6fafe49",
  1152 => x"87c4c187",
  1153 => x"91cb4974",
  1154 => x"81dee4c1",
  1155 => x"79dfc0c1",
  1156 => x"97dee3c2",
  1157 => x"87d802bf",
  1158 => x"91de4974",
  1159 => x"e8c284c1",
  1160 => x"83714bec",
  1161 => x"4adee3c2",
  1162 => x"f9fe49dd",
  1163 => x"87d887f9",
  1164 => x"93de4b74",
  1165 => x"83ece8c2",
  1166 => x"c049a3cb",
  1167 => x"7384c151",
  1168 => x"49cb4a6e",
  1169 => x"87dff9fe",
  1170 => x"c14866c4",
  1171 => x"58a6c880",
  1172 => x"c003acc7",
  1173 => x"056e87c5",
  1174 => x"7487e4fc",
  1175 => x"f48ef448",
  1176 => x"731e87f6",
  1177 => x"494b711e",
  1178 => x"e4c191cb",
  1179 => x"a1c881de",
  1180 => x"cae4c14a",
  1181 => x"c9501248",
  1182 => x"f9c04aa1",
  1183 => x"501248c0",
  1184 => x"e4c181ca",
  1185 => x"501148cb",
  1186 => x"97cbe4c1",
  1187 => x"c01e49bf",
  1188 => x"87cbf549",
  1189 => x"48c0e8c2",
  1190 => x"49c178de",
  1191 => x"2687efd5",
  1192 => x"0e87f9f3",
  1193 => x"5d5c5b5e",
  1194 => x"7186f40e",
  1195 => x"91cb494d",
  1196 => x"81dee4c1",
  1197 => x"ca4aa1c8",
  1198 => x"a6c47ea1",
  1199 => x"c8ecc248",
  1200 => x"976e78bf",
  1201 => x"66c44bbf",
  1202 => x"122c734c",
  1203 => x"58a6cc48",
  1204 => x"84c19c70",
  1205 => x"699781c9",
  1206 => x"04acb749",
  1207 => x"4cc087c2",
  1208 => x"4abf976e",
  1209 => x"724966c8",
  1210 => x"c4b9ff31",
  1211 => x"48749966",
  1212 => x"4a703072",
  1213 => x"c2b07148",
  1214 => x"c058ccec",
  1215 => x"c087d8e5",
  1216 => x"87cad449",
  1217 => x"f7c04975",
  1218 => x"8ef487cd",
  1219 => x"1e87c9f2",
  1220 => x"4b711e73",
  1221 => x"87cbfe49",
  1222 => x"c6fe4973",
  1223 => x"87fcf187",
  1224 => x"711e731e",
  1225 => x"4aa3c64b",
  1226 => x"c187db02",
  1227 => x"87d6028a",
  1228 => x"dac1028a",
  1229 => x"c0028a87",
  1230 => x"028a87fc",
  1231 => x"8a87e1c0",
  1232 => x"c187cb02",
  1233 => x"49c787db",
  1234 => x"c187c7f6",
  1235 => x"e8c287de",
  1236 => x"c102bfd8",
  1237 => x"c14887cb",
  1238 => x"dce8c288",
  1239 => x"87c1c158",
  1240 => x"bfdce8c2",
  1241 => x"87f9c002",
  1242 => x"bfd8e8c2",
  1243 => x"c280c148",
  1244 => x"c058dce8",
  1245 => x"e8c287eb",
  1246 => x"c649bfd8",
  1247 => x"dce8c289",
  1248 => x"a9b7c059",
  1249 => x"c287da03",
  1250 => x"c048d8e8",
  1251 => x"c287d278",
  1252 => x"02bfdce8",
  1253 => x"e8c287cb",
  1254 => x"c648bfd8",
  1255 => x"dce8c280",
  1256 => x"d149c058",
  1257 => x"497387e8",
  1258 => x"87ebf4c0",
  1259 => x"0e87edef",
  1260 => x"5d5c5b5e",
  1261 => x"86d4ff0e",
  1262 => x"c859a6dc",
  1263 => x"78c048a6",
  1264 => x"c0c180c4",
  1265 => x"80c47866",
  1266 => x"80c478c1",
  1267 => x"e8c278c1",
  1268 => x"78c148dc",
  1269 => x"bfc0e8c2",
  1270 => x"05a8de48",
  1271 => x"f8f487c9",
  1272 => x"58a6cc87",
  1273 => x"e387e6cf",
  1274 => x"fbe387d9",
  1275 => x"87c8e387",
  1276 => x"fbc04c70",
  1277 => x"fbc102ac",
  1278 => x"0566d887",
  1279 => x"c087edc1",
  1280 => x"c44a66fc",
  1281 => x"727e6a82",
  1282 => x"c2e0c11e",
  1283 => x"4966c448",
  1284 => x"204aa1c8",
  1285 => x"05aa7141",
  1286 => x"511087f9",
  1287 => x"fcc04a26",
  1288 => x"c9c14866",
  1289 => x"496a78e2",
  1290 => x"517481c7",
  1291 => x"4966fcc0",
  1292 => x"51c181c8",
  1293 => x"4966fcc0",
  1294 => x"51c081c9",
  1295 => x"4966fcc0",
  1296 => x"51c081ca",
  1297 => x"1ed81ec1",
  1298 => x"81c8496a",
  1299 => x"c887ede2",
  1300 => x"66c0c186",
  1301 => x"01a8c048",
  1302 => x"a6c887c7",
  1303 => x"ce78c148",
  1304 => x"66c0c187",
  1305 => x"d088c148",
  1306 => x"87c358a6",
  1307 => x"d087f9e1",
  1308 => x"78c248a6",
  1309 => x"cd029c74",
  1310 => x"66c887cf",
  1311 => x"66c4c148",
  1312 => x"c4cd03a8",
  1313 => x"48a6dc87",
  1314 => x"80e878c0",
  1315 => x"e7e078c0",
  1316 => x"c14c7087",
  1317 => x"c205acd0",
  1318 => x"66c487d7",
  1319 => x"87cbe37e",
  1320 => x"e058a6c8",
  1321 => x"4c7087d2",
  1322 => x"05acecc0",
  1323 => x"c887edc1",
  1324 => x"91cb4966",
  1325 => x"8166fcc0",
  1326 => x"6a4aa1c4",
  1327 => x"4aa1c84d",
  1328 => x"c15266c4",
  1329 => x"ff79d2c3",
  1330 => x"7087eddf",
  1331 => x"d9029c4c",
  1332 => x"acfbc087",
  1333 => x"7487d302",
  1334 => x"dbdfff55",
  1335 => x"9c4c7087",
  1336 => x"c087c702",
  1337 => x"ff05acfb",
  1338 => x"e0c087ed",
  1339 => x"55c1c255",
  1340 => x"d87d97c0",
  1341 => x"a86e4866",
  1342 => x"c887db05",
  1343 => x"66cc4866",
  1344 => x"87ca04a8",
  1345 => x"c14866c8",
  1346 => x"58a6cc80",
  1347 => x"66cc87c8",
  1348 => x"d088c148",
  1349 => x"deff58a6",
  1350 => x"4c7087de",
  1351 => x"05acd0c1",
  1352 => x"66d487c8",
  1353 => x"d880c148",
  1354 => x"d0c158a6",
  1355 => x"e9fd02ac",
  1356 => x"4866c487",
  1357 => x"05a866d8",
  1358 => x"c087e0c9",
  1359 => x"c048a6e0",
  1360 => x"c0487478",
  1361 => x"7e7088fb",
  1362 => x"c9029848",
  1363 => x"cb4887e2",
  1364 => x"487e7088",
  1365 => x"cdc10298",
  1366 => x"88c94887",
  1367 => x"98487e70",
  1368 => x"87fec302",
  1369 => x"7088c448",
  1370 => x"0298487e",
  1371 => x"c14887ce",
  1372 => x"487e7088",
  1373 => x"e9c30298",
  1374 => x"87d6c887",
  1375 => x"c048a6dc",
  1376 => x"dcff78f0",
  1377 => x"4c7087f2",
  1378 => x"02acecc0",
  1379 => x"c087c4c0",
  1380 => x"c05ca6e0",
  1381 => x"cd02acec",
  1382 => x"dbdcff87",
  1383 => x"c04c7087",
  1384 => x"ff05acec",
  1385 => x"ecc087f3",
  1386 => x"c4c002ac",
  1387 => x"c7dcff87",
  1388 => x"ca1ec087",
  1389 => x"4966d01e",
  1390 => x"c4c191cb",
  1391 => x"80714866",
  1392 => x"c858a6cc",
  1393 => x"80c44866",
  1394 => x"cc58a6d0",
  1395 => x"ff49bf66",
  1396 => x"c187e9dc",
  1397 => x"d41ede1e",
  1398 => x"ff49bf66",
  1399 => x"d087dddc",
  1400 => x"48497086",
  1401 => x"c08808c0",
  1402 => x"c058a6e8",
  1403 => x"eec006a8",
  1404 => x"66e4c087",
  1405 => x"03a8dd48",
  1406 => x"c487e4c0",
  1407 => x"c049bf66",
  1408 => x"c08166e4",
  1409 => x"e4c051e0",
  1410 => x"81c14966",
  1411 => x"81bf66c4",
  1412 => x"c051c1c2",
  1413 => x"c24966e4",
  1414 => x"bf66c481",
  1415 => x"6e51c081",
  1416 => x"e2c9c148",
  1417 => x"c8496e78",
  1418 => x"5166d081",
  1419 => x"81c9496e",
  1420 => x"6e5166d4",
  1421 => x"dc81ca49",
  1422 => x"66d05166",
  1423 => x"d480c148",
  1424 => x"66c858a6",
  1425 => x"a866cc48",
  1426 => x"87cbc004",
  1427 => x"c14866c8",
  1428 => x"58a6cc80",
  1429 => x"cc87d9c5",
  1430 => x"88c14866",
  1431 => x"c558a6d0",
  1432 => x"dcff87ce",
  1433 => x"e8c087c5",
  1434 => x"dbff58a6",
  1435 => x"e0c087fd",
  1436 => x"ecc058a6",
  1437 => x"cac005a8",
  1438 => x"48a6dc87",
  1439 => x"7866e4c0",
  1440 => x"ff87c4c0",
  1441 => x"c887f1d8",
  1442 => x"91cb4966",
  1443 => x"4866fcc0",
  1444 => x"7e708071",
  1445 => x"6e82c84a",
  1446 => x"c081ca49",
  1447 => x"dc5166e4",
  1448 => x"81c14966",
  1449 => x"8966e4c0",
  1450 => x"307148c1",
  1451 => x"89c14970",
  1452 => x"c27a9771",
  1453 => x"49bfc8ec",
  1454 => x"2966e4c0",
  1455 => x"484a6a97",
  1456 => x"ecc09871",
  1457 => x"496e58a6",
  1458 => x"4d6981c4",
  1459 => x"c44866d8",
  1460 => x"c002a866",
  1461 => x"a6c487c8",
  1462 => x"c078c048",
  1463 => x"a6c487c5",
  1464 => x"c478c148",
  1465 => x"e0c01e66",
  1466 => x"ff49751e",
  1467 => x"c887cdd8",
  1468 => x"c04c7086",
  1469 => x"c106acb7",
  1470 => x"857487d4",
  1471 => x"7449e0c0",
  1472 => x"c14b7589",
  1473 => x"714acbe0",
  1474 => x"87dbe6fe",
  1475 => x"e0c085c2",
  1476 => x"80c14866",
  1477 => x"58a6e4c0",
  1478 => x"4966e8c0",
  1479 => x"a97081c1",
  1480 => x"87c8c002",
  1481 => x"c048a6c4",
  1482 => x"87c5c078",
  1483 => x"c148a6c4",
  1484 => x"1e66c478",
  1485 => x"c049a4c2",
  1486 => x"887148e0",
  1487 => x"751e4970",
  1488 => x"f7d6ff49",
  1489 => x"c086c887",
  1490 => x"ff01a8b7",
  1491 => x"e0c087c0",
  1492 => x"d1c00266",
  1493 => x"c9496e87",
  1494 => x"66e0c081",
  1495 => x"c1486e51",
  1496 => x"c078e3ca",
  1497 => x"496e87cc",
  1498 => x"51c281c9",
  1499 => x"ccc1486e",
  1500 => x"66c878cf",
  1501 => x"a866cc48",
  1502 => x"87cbc004",
  1503 => x"c14866c8",
  1504 => x"58a6cc80",
  1505 => x"cc87e9c0",
  1506 => x"88c14866",
  1507 => x"c058a6d0",
  1508 => x"d5ff87de",
  1509 => x"4c7087d2",
  1510 => x"c187d5c0",
  1511 => x"c005acc6",
  1512 => x"66d087c8",
  1513 => x"d480c148",
  1514 => x"d4ff58a6",
  1515 => x"4c7087fa",
  1516 => x"c14866d4",
  1517 => x"58a6d880",
  1518 => x"c0029c74",
  1519 => x"66c887cb",
  1520 => x"66c4c148",
  1521 => x"fcf204a8",
  1522 => x"d2d4ff87",
  1523 => x"4866c887",
  1524 => x"c003a8c7",
  1525 => x"e8c287e5",
  1526 => x"78c048dc",
  1527 => x"cb4966c8",
  1528 => x"66fcc091",
  1529 => x"4aa1c481",
  1530 => x"52c04a6a",
  1531 => x"4866c879",
  1532 => x"a6cc80c1",
  1533 => x"04a8c758",
  1534 => x"ff87dbff",
  1535 => x"deff8ed4",
  1536 => x"6f4c87d6",
  1537 => x"2a206461",
  1538 => x"3a00202e",
  1539 => x"731e0020",
  1540 => x"9b4b711e",
  1541 => x"c287c602",
  1542 => x"c048d8e8",
  1543 => x"c21ec778",
  1544 => x"1ebfd8e8",
  1545 => x"1edee4c1",
  1546 => x"bfc0e8c2",
  1547 => x"87ffed49",
  1548 => x"e8c286cc",
  1549 => x"e249bfc0",
  1550 => x"9b7387f7",
  1551 => x"c187c802",
  1552 => x"c049dee4",
  1553 => x"ff87e2e3",
  1554 => x"1e87d1dd",
  1555 => x"4bc01e73",
  1556 => x"48cae4c1",
  1557 => x"e6c150c0",
  1558 => x"ff49bfc1",
  1559 => x"7087e2d7",
  1560 => x"87c40598",
  1561 => x"4beee1c1",
  1562 => x"dcff4873",
  1563 => x"4f5287ee",
  1564 => x"6f6c204d",
  1565 => x"6e696461",
  1566 => x"61662067",
  1567 => x"64656c69",
  1568 => x"e3c71e00",
  1569 => x"fe49c187",
  1570 => x"e9fe87c4",
  1571 => x"987087c9",
  1572 => x"fe87cd02",
  1573 => x"7087c3f2",
  1574 => x"87c40298",
  1575 => x"87c24ac1",
  1576 => x"9a724ac0",
  1577 => x"c087ce05",
  1578 => x"d1e3c11e",
  1579 => x"eeeec049",
  1580 => x"fe86c487",
  1581 => x"c11ec087",
  1582 => x"c049dce3",
  1583 => x"c087e0ee",
  1584 => x"87c7fe1e",
  1585 => x"eec04970",
  1586 => x"dac387d5",
  1587 => x"268ef887",
  1588 => x"2044534f",
  1589 => x"6c696166",
  1590 => x"002e6465",
  1591 => x"746f6f42",
  1592 => x"2e676e69",
  1593 => x"1e002e2e",
  1594 => x"87fae5c0",
  1595 => x"87e9f1c0",
  1596 => x"4f2687f6",
  1597 => x"d8e8c21e",
  1598 => x"c278c048",
  1599 => x"c048c0e8",
  1600 => x"87fdfd78",
  1601 => x"48c087e1",
  1602 => x"00004f26",
  1603 => x"00000001",
  1604 => x"78452080",
  1605 => x"80007469",
  1606 => x"63614220",
  1607 => x"101f006b",
  1608 => x"2a2c0000",
  1609 => x"00000000",
  1610 => x"00101f00",
  1611 => x"002a4a00",
  1612 => x"00000000",
  1613 => x"0000101f",
  1614 => x"00002a68",
  1615 => x"1f000000",
  1616 => x"86000010",
  1617 => x"0000002a",
  1618 => x"101f0000",
  1619 => x"2aa40000",
  1620 => x"00000000",
  1621 => x"00101f00",
  1622 => x"002ac200",
  1623 => x"00000000",
  1624 => x"0000101f",
  1625 => x"00002ae0",
  1626 => x"d2000000",
  1627 => x"00000010",
  1628 => x"00000000",
  1629 => x"13200000",
  1630 => x"00000000",
  1631 => x"00000000",
  1632 => x"00198500",
  1633 => x"39495400",
  1634 => x"20413439",
  1635 => x"4d4f5220",
  1636 => x"f0fe1e00",
  1637 => x"cd78c048",
  1638 => x"26097909",
  1639 => x"fe1e1e4f",
  1640 => x"487ebff0",
  1641 => x"1e4f2626",
  1642 => x"c148f0fe",
  1643 => x"1e4f2678",
  1644 => x"c048f0fe",
  1645 => x"1e4f2678",
  1646 => x"52c04a71",
  1647 => x"0e4f2652",
  1648 => x"5d5c5b5e",
  1649 => x"7186f40e",
  1650 => x"7e6d974d",
  1651 => x"974ca5c1",
  1652 => x"a6c8486c",
  1653 => x"c4486e58",
  1654 => x"c505a866",
  1655 => x"c048ff87",
  1656 => x"caff87e6",
  1657 => x"49a5c287",
  1658 => x"714b6c97",
  1659 => x"6b974ba3",
  1660 => x"7e6c974b",
  1661 => x"80c1486e",
  1662 => x"c758a6c8",
  1663 => x"58a6cc98",
  1664 => x"fe7c9770",
  1665 => x"487387e1",
  1666 => x"4d268ef4",
  1667 => x"4b264c26",
  1668 => x"5e0e4f26",
  1669 => x"f40e5c5b",
  1670 => x"d84c7186",
  1671 => x"ffc34a66",
  1672 => x"4ba4c29a",
  1673 => x"73496c97",
  1674 => x"517249a1",
  1675 => x"6e7e6c97",
  1676 => x"c880c148",
  1677 => x"98c758a6",
  1678 => x"7058a6cc",
  1679 => x"ff8ef454",
  1680 => x"1e1e87ca",
  1681 => x"e087e8fd",
  1682 => x"c0494abf",
  1683 => x"0299c0e0",
  1684 => x"1e7287cb",
  1685 => x"49feebc2",
  1686 => x"c487f7fe",
  1687 => x"87fdfc86",
  1688 => x"c2fd7e70",
  1689 => x"4f262687",
  1690 => x"feebc21e",
  1691 => x"87c7fd49",
  1692 => x"49c2e9c1",
  1693 => x"c387dafc",
  1694 => x"4f2687f7",
  1695 => x"5c5b5e0e",
  1696 => x"4d710e5d",
  1697 => x"49feebc2",
  1698 => x"7087f4fc",
  1699 => x"abb7c04b",
  1700 => x"87c2c304",
  1701 => x"05abf0c3",
  1702 => x"edc187c9",
  1703 => x"78c148e0",
  1704 => x"c387e3c2",
  1705 => x"c905abe0",
  1706 => x"e4edc187",
  1707 => x"c278c148",
  1708 => x"edc187d4",
  1709 => x"c602bfe4",
  1710 => x"a3c0c287",
  1711 => x"7387c24c",
  1712 => x"e0edc14c",
  1713 => x"e0c002bf",
  1714 => x"c4497487",
  1715 => x"c19129b7",
  1716 => x"7481c0ef",
  1717 => x"c29acf4a",
  1718 => x"7248c192",
  1719 => x"ff4a7030",
  1720 => x"694872ba",
  1721 => x"db797098",
  1722 => x"c4497487",
  1723 => x"c19129b7",
  1724 => x"7481c0ef",
  1725 => x"c29acf4a",
  1726 => x"7248c392",
  1727 => x"484a7030",
  1728 => x"7970b069",
  1729 => x"c0059d75",
  1730 => x"d0ff87f0",
  1731 => x"78e1c848",
  1732 => x"c548d4ff",
  1733 => x"e4edc178",
  1734 => x"87c302bf",
  1735 => x"c178e0c3",
  1736 => x"02bfe0ed",
  1737 => x"d4ff87c6",
  1738 => x"78f0c348",
  1739 => x"7b0bd4ff",
  1740 => x"48d0ff0b",
  1741 => x"c078e1c8",
  1742 => x"edc178e0",
  1743 => x"78c048e4",
  1744 => x"48e0edc1",
  1745 => x"ebc278c0",
  1746 => x"f2f949fe",
  1747 => x"c04b7087",
  1748 => x"fc03abb7",
  1749 => x"48c087fe",
  1750 => x"4c264d26",
  1751 => x"4f264b26",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"494a711e",
  1755 => x"2687cdfc",
  1756 => x"4ac01e4f",
  1757 => x"91c44972",
  1758 => x"81c0efc1",
  1759 => x"82c179c0",
  1760 => x"04aab7d0",
  1761 => x"4f2687ee",
  1762 => x"5c5b5e0e",
  1763 => x"4d710e5d",
  1764 => x"7587dcf8",
  1765 => x"2ab7c44a",
  1766 => x"c0efc192",
  1767 => x"cf4c7582",
  1768 => x"6a94c29c",
  1769 => x"2b744b49",
  1770 => x"48c29bc3",
  1771 => x"4c703074",
  1772 => x"4874bcff",
  1773 => x"7a709871",
  1774 => x"7387ecf7",
  1775 => x"87d8fe48",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"48d0ff1e",
  1793 => x"7178e1c8",
  1794 => x"08d4ff48",
  1795 => x"1e4f2678",
  1796 => x"c848d0ff",
  1797 => x"487178e1",
  1798 => x"7808d4ff",
  1799 => x"ff4866c4",
  1800 => x"267808d4",
  1801 => x"4a711e4f",
  1802 => x"1e4966c4",
  1803 => x"deff4972",
  1804 => x"48d0ff87",
  1805 => x"2678e0c0",
  1806 => x"731e4f26",
  1807 => x"c84b711e",
  1808 => x"731e4966",
  1809 => x"a2e0c14a",
  1810 => x"87d9ff49",
  1811 => x"2687c426",
  1812 => x"264c264d",
  1813 => x"1e4f264b",
  1814 => x"c34ad4ff",
  1815 => x"d0ff7aff",
  1816 => x"78e1c048",
  1817 => x"ecc27ade",
  1818 => x"497abfc8",
  1819 => x"7028c848",
  1820 => x"d048717a",
  1821 => x"717a7028",
  1822 => x"7028d848",
  1823 => x"48d0ff7a",
  1824 => x"2678e0c0",
  1825 => x"d0ff1e4f",
  1826 => x"78c9c848",
  1827 => x"d4ff4871",
  1828 => x"4f267808",
  1829 => x"494a711e",
  1830 => x"d0ff87eb",
  1831 => x"2678c848",
  1832 => x"1e731e4f",
  1833 => x"ecc24b71",
  1834 => x"c302bfd8",
  1835 => x"87ebc287",
  1836 => x"c848d0ff",
  1837 => x"487378c9",
  1838 => x"ffb0e0c0",
  1839 => x"c27808d4",
  1840 => x"c048ccec",
  1841 => x"0266c878",
  1842 => x"ffc387c5",
  1843 => x"c087c249",
  1844 => x"d4ecc249",
  1845 => x"0266cc59",
  1846 => x"d5c587c6",
  1847 => x"87c44ad5",
  1848 => x"4affffcf",
  1849 => x"5ad8ecc2",
  1850 => x"48d8ecc2",
  1851 => x"87c478c1",
  1852 => x"4c264d26",
  1853 => x"4f264b26",
  1854 => x"5c5b5e0e",
  1855 => x"4a710e5d",
  1856 => x"bfd4ecc2",
  1857 => x"029a724c",
  1858 => x"c84987cb",
  1859 => x"d7f2c191",
  1860 => x"c483714b",
  1861 => x"d7f6c187",
  1862 => x"134dc04b",
  1863 => x"c2997449",
  1864 => x"48bfd0ec",
  1865 => x"d4ffb871",
  1866 => x"b7c17808",
  1867 => x"b7c8852c",
  1868 => x"87e704ad",
  1869 => x"bfccecc2",
  1870 => x"c280c848",
  1871 => x"fe58d0ec",
  1872 => x"731e87ee",
  1873 => x"134b711e",
  1874 => x"cb029a4a",
  1875 => x"fe497287",
  1876 => x"4a1387e6",
  1877 => x"87f5059a",
  1878 => x"1e87d9fe",
  1879 => x"bfccecc2",
  1880 => x"ccecc249",
  1881 => x"78a1c148",
  1882 => x"a9b7c0c4",
  1883 => x"ff87db03",
  1884 => x"ecc248d4",
  1885 => x"c278bfd0",
  1886 => x"49bfccec",
  1887 => x"48ccecc2",
  1888 => x"c478a1c1",
  1889 => x"04a9b7c0",
  1890 => x"d0ff87e5",
  1891 => x"c278c848",
  1892 => x"c048d8ec",
  1893 => x"004f2678",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"5f5f0000",
  1897 => x"00000000",
  1898 => x"03000303",
  1899 => x"14000003",
  1900 => x"7f147f7f",
  1901 => x"0000147f",
  1902 => x"6b6b2e24",
  1903 => x"4c00123a",
  1904 => x"6c18366a",
  1905 => x"30003256",
  1906 => x"77594f7e",
  1907 => x"0040683a",
  1908 => x"03070400",
  1909 => x"00000000",
  1910 => x"633e1c00",
  1911 => x"00000041",
  1912 => x"3e634100",
  1913 => x"0800001c",
  1914 => x"1c1c3e2a",
  1915 => x"00082a3e",
  1916 => x"3e3e0808",
  1917 => x"00000808",
  1918 => x"60e08000",
  1919 => x"00000000",
  1920 => x"08080808",
  1921 => x"00000808",
  1922 => x"60600000",
  1923 => x"40000000",
  1924 => x"0c183060",
  1925 => x"00010306",
  1926 => x"4d597f3e",
  1927 => x"00003e7f",
  1928 => x"7f7f0604",
  1929 => x"00000000",
  1930 => x"59716342",
  1931 => x"0000464f",
  1932 => x"49496322",
  1933 => x"1800367f",
  1934 => x"7f13161c",
  1935 => x"0000107f",
  1936 => x"45456727",
  1937 => x"0000397d",
  1938 => x"494b7e3c",
  1939 => x"00003079",
  1940 => x"79710101",
  1941 => x"0000070f",
  1942 => x"49497f36",
  1943 => x"0000367f",
  1944 => x"69494f06",
  1945 => x"00001e3f",
  1946 => x"66660000",
  1947 => x"00000000",
  1948 => x"66e68000",
  1949 => x"00000000",
  1950 => x"14140808",
  1951 => x"00002222",
  1952 => x"14141414",
  1953 => x"00001414",
  1954 => x"14142222",
  1955 => x"00000808",
  1956 => x"59510302",
  1957 => x"3e00060f",
  1958 => x"555d417f",
  1959 => x"00001e1f",
  1960 => x"09097f7e",
  1961 => x"00007e7f",
  1962 => x"49497f7f",
  1963 => x"0000367f",
  1964 => x"41633e1c",
  1965 => x"00004141",
  1966 => x"63417f7f",
  1967 => x"00001c3e",
  1968 => x"49497f7f",
  1969 => x"00004141",
  1970 => x"09097f7f",
  1971 => x"00000101",
  1972 => x"49417f3e",
  1973 => x"00007a7b",
  1974 => x"08087f7f",
  1975 => x"00007f7f",
  1976 => x"7f7f4100",
  1977 => x"00000041",
  1978 => x"40406020",
  1979 => x"7f003f7f",
  1980 => x"361c087f",
  1981 => x"00004163",
  1982 => x"40407f7f",
  1983 => x"7f004040",
  1984 => x"060c067f",
  1985 => x"7f007f7f",
  1986 => x"180c067f",
  1987 => x"00007f7f",
  1988 => x"41417f3e",
  1989 => x"00003e7f",
  1990 => x"09097f7f",
  1991 => x"3e00060f",
  1992 => x"7f61417f",
  1993 => x"0000407e",
  1994 => x"19097f7f",
  1995 => x"0000667f",
  1996 => x"594d6f26",
  1997 => x"0000327b",
  1998 => x"7f7f0101",
  1999 => x"00000101",
  2000 => x"40407f3f",
  2001 => x"00003f7f",
  2002 => x"70703f0f",
  2003 => x"7f000f3f",
  2004 => x"3018307f",
  2005 => x"41007f7f",
  2006 => x"1c1c3663",
  2007 => x"01416336",
  2008 => x"7c7c0603",
  2009 => x"61010306",
  2010 => x"474d5971",
  2011 => x"00004143",
  2012 => x"417f7f00",
  2013 => x"01000041",
  2014 => x"180c0603",
  2015 => x"00406030",
  2016 => x"7f414100",
  2017 => x"0800007f",
  2018 => x"0603060c",
  2019 => x"8000080c",
  2020 => x"80808080",
  2021 => x"00008080",
  2022 => x"07030000",
  2023 => x"00000004",
  2024 => x"54547420",
  2025 => x"0000787c",
  2026 => x"44447f7f",
  2027 => x"0000387c",
  2028 => x"44447c38",
  2029 => x"00000044",
  2030 => x"44447c38",
  2031 => x"00007f7f",
  2032 => x"54547c38",
  2033 => x"0000185c",
  2034 => x"057f7e04",
  2035 => x"00000005",
  2036 => x"a4a4bc18",
  2037 => x"00007cfc",
  2038 => x"04047f7f",
  2039 => x"0000787c",
  2040 => x"7d3d0000",
  2041 => x"00000040",
  2042 => x"fd808080",
  2043 => x"0000007d",
  2044 => x"38107f7f",
  2045 => x"0000446c",
  2046 => x"7f3f0000",
  2047 => x"7c000040",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
