library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0c180c7c",
     1 => x"0000787c",
     2 => x"04047c7c",
     3 => x"0000787c",
     4 => x"44447c38",
     5 => x"0000387c",
     6 => x"2424fcfc",
     7 => x"0000183c",
     8 => x"24243c18",
     9 => x"0000fcfc",
    10 => x"04047c7c",
    11 => x"0000080c",
    12 => x"54545c48",
    13 => x"00002074",
    14 => x"447f3f04",
    15 => x"00000044",
    16 => x"40407c3c",
    17 => x"00007c7c",
    18 => x"60603c1c",
    19 => x"3c001c3c",
    20 => x"6030607c",
    21 => x"44003c7c",
    22 => x"3810386c",
    23 => x"0000446c",
    24 => x"60e0bc1c",
    25 => x"00001c3c",
    26 => x"5c746444",
    27 => x"0000444c",
    28 => x"773e0808",
    29 => x"00004141",
    30 => x"7f7f0000",
    31 => x"00000000",
    32 => x"3e774141",
    33 => x"02000808",
    34 => x"02030101",
    35 => x"7f000102",
    36 => x"7f7f7f7f",
    37 => x"08007f7f",
    38 => x"3e1c1c08",
    39 => x"7f7f7f3e",
    40 => x"1c3e3e7f",
    41 => x"0008081c",
    42 => x"7c7c1810",
    43 => x"00001018",
    44 => x"7c7c3010",
    45 => x"10001030",
    46 => x"78606030",
    47 => x"4200061e",
    48 => x"3c183c66",
    49 => x"78004266",
    50 => x"c6c26a38",
    51 => x"6000386c",
    52 => x"00600000",
    53 => x"0e006000",
    54 => x"5d5c5b5e",
    55 => x"4c711e0e",
    56 => x"bfe9ecc2",
    57 => x"c04bc04d",
    58 => x"02ab741e",
    59 => x"a6c487c7",
    60 => x"c578c048",
    61 => x"48a6c487",
    62 => x"66c478c1",
    63 => x"ee49731e",
    64 => x"86c887df",
    65 => x"ef49e0c0",
    66 => x"a5c487ee",
    67 => x"f0496a4a",
    68 => x"c6f187f0",
    69 => x"c185cb87",
    70 => x"abb7c883",
    71 => x"87c7ff04",
    72 => x"264d2626",
    73 => x"264b264c",
    74 => x"4a711e4f",
    75 => x"5aedecc2",
    76 => x"48edecc2",
    77 => x"fe4978c7",
    78 => x"4f2687dd",
    79 => x"711e731e",
    80 => x"aab7c04a",
    81 => x"c287d303",
    82 => x"05bff8d2",
    83 => x"4bc187c4",
    84 => x"4bc087c2",
    85 => x"5bfcd2c2",
    86 => x"d2c287c4",
    87 => x"d2c25afc",
    88 => x"c14abff8",
    89 => x"a2c0c19a",
    90 => x"87e8ec49",
    91 => x"d2c248fc",
    92 => x"fe78bff8",
    93 => x"711e87ef",
    94 => x"1e66c44a",
    95 => x"f9ea4972",
    96 => x"4f262687",
    97 => x"48d4ff1e",
    98 => x"ff78ffc3",
    99 => x"e1c048d0",
   100 => x"48d4ff78",
   101 => x"487178c1",
   102 => x"d4ff30c4",
   103 => x"d0ff7808",
   104 => x"78e0c048",
   105 => x"c21e4f26",
   106 => x"49bff8d2",
   107 => x"c287f9e6",
   108 => x"e848e1ec",
   109 => x"ecc278bf",
   110 => x"bfec48dd",
   111 => x"e1ecc278",
   112 => x"c3494abf",
   113 => x"b7c899ff",
   114 => x"7148722a",
   115 => x"e9ecc2b0",
   116 => x"0e4f2658",
   117 => x"5d5c5b5e",
   118 => x"ff4b710e",
   119 => x"ecc287c8",
   120 => x"50c048dc",
   121 => x"dfe64973",
   122 => x"4c497087",
   123 => x"eecb9cc2",
   124 => x"87cccb49",
   125 => x"ecc24d70",
   126 => x"05bf97dc",
   127 => x"d087e2c1",
   128 => x"ecc24966",
   129 => x"0599bfe5",
   130 => x"66d487d6",
   131 => x"ddecc249",
   132 => x"cb0599bf",
   133 => x"e5497387",
   134 => x"987087ee",
   135 => x"87c1c102",
   136 => x"c1fe4cc1",
   137 => x"ca497587",
   138 => x"987087e2",
   139 => x"c287c602",
   140 => x"c148dcec",
   141 => x"dcecc250",
   142 => x"c005bf97",
   143 => x"ecc287e3",
   144 => x"d049bfe5",
   145 => x"ff059966",
   146 => x"ecc287d6",
   147 => x"d449bfdd",
   148 => x"ff059966",
   149 => x"497387ca",
   150 => x"7087ede4",
   151 => x"fffe0598",
   152 => x"fa487487",
   153 => x"5e0e87fb",
   154 => x"0e5d5c5b",
   155 => x"4dc086f8",
   156 => x"7ebfec4c",
   157 => x"c248a6c4",
   158 => x"78bfe9ec",
   159 => x"1ec01ec1",
   160 => x"cefd49c7",
   161 => x"7086c887",
   162 => x"87cd0298",
   163 => x"ebfa49ff",
   164 => x"49dac187",
   165 => x"c187f1e3",
   166 => x"dcecc24d",
   167 => x"cf02bf97",
   168 => x"f0d2c287",
   169 => x"b9c149bf",
   170 => x"59f4d2c2",
   171 => x"87d4fb71",
   172 => x"bfe1ecc2",
   173 => x"f8d2c24b",
   174 => x"e9c005bf",
   175 => x"49fdc387",
   176 => x"c387c5e3",
   177 => x"ffe249fa",
   178 => x"c3497387",
   179 => x"1e7199ff",
   180 => x"e1fa49c0",
   181 => x"c8497387",
   182 => x"1e7129b7",
   183 => x"d5fa49c1",
   184 => x"c586c887",
   185 => x"ecc287f4",
   186 => x"9b4bbfe5",
   187 => x"c287dd02",
   188 => x"49bff4d2",
   189 => x"7087d5c7",
   190 => x"87c40598",
   191 => x"87d24bc0",
   192 => x"c649e0c2",
   193 => x"d2c287fa",
   194 => x"87c658f8",
   195 => x"48f4d2c2",
   196 => x"497378c0",
   197 => x"cd0599c2",
   198 => x"49ebc387",
   199 => x"7087e9e1",
   200 => x"0299c249",
   201 => x"4cfb87c2",
   202 => x"99c14973",
   203 => x"c387cd05",
   204 => x"d3e149f4",
   205 => x"c2497087",
   206 => x"87c20299",
   207 => x"49734cfa",
   208 => x"cd0599c8",
   209 => x"49f5c387",
   210 => x"7087fde0",
   211 => x"0299c249",
   212 => x"ecc287d5",
   213 => x"ca02bfed",
   214 => x"88c14887",
   215 => x"58f1ecc2",
   216 => x"ff87c2c0",
   217 => x"734dc14c",
   218 => x"0599c449",
   219 => x"f2c387cd",
   220 => x"87d4e049",
   221 => x"99c24970",
   222 => x"c287dc02",
   223 => x"7ebfedec",
   224 => x"a8b7c748",
   225 => x"87cbc003",
   226 => x"80c1486e",
   227 => x"58f1ecc2",
   228 => x"fe87c2c0",
   229 => x"c34dc14c",
   230 => x"dfff49fd",
   231 => x"497087ea",
   232 => x"d50299c2",
   233 => x"edecc287",
   234 => x"c9c002bf",
   235 => x"edecc287",
   236 => x"c078c048",
   237 => x"4cfd87c2",
   238 => x"fac34dc1",
   239 => x"c7dfff49",
   240 => x"c2497087",
   241 => x"d9c00299",
   242 => x"edecc287",
   243 => x"b7c748bf",
   244 => x"c9c003a8",
   245 => x"edecc287",
   246 => x"c078c748",
   247 => x"4cfc87c2",
   248 => x"b7c04dc1",
   249 => x"d3c003ac",
   250 => x"4866c487",
   251 => x"7080d8c1",
   252 => x"02bf6e7e",
   253 => x"4b87c5c0",
   254 => x"0f734974",
   255 => x"f0c31ec0",
   256 => x"49dac11e",
   257 => x"c887ccf7",
   258 => x"02987086",
   259 => x"c287d8c0",
   260 => x"7ebfedec",
   261 => x"91cb496e",
   262 => x"714a66c4",
   263 => x"c0026a82",
   264 => x"6e4b87c5",
   265 => x"750f7349",
   266 => x"c8c0029d",
   267 => x"edecc287",
   268 => x"e2f249bf",
   269 => x"fcd2c287",
   270 => x"ddc002bf",
   271 => x"cbc24987",
   272 => x"02987087",
   273 => x"c287d3c0",
   274 => x"49bfedec",
   275 => x"c087c8f2",
   276 => x"87e8f349",
   277 => x"48fcd2c2",
   278 => x"8ef878c0",
   279 => x"0e87c2f3",
   280 => x"5d5c5b5e",
   281 => x"4c711e0e",
   282 => x"bfe9ecc2",
   283 => x"a1cdc149",
   284 => x"81d1c14d",
   285 => x"9c747e69",
   286 => x"c487cf02",
   287 => x"7b744ba5",
   288 => x"bfe9ecc2",
   289 => x"87e1f249",
   290 => x"9c747b6e",
   291 => x"c087c405",
   292 => x"c187c24b",
   293 => x"f249734b",
   294 => x"66d487e2",
   295 => x"4987c702",
   296 => x"4a7087de",
   297 => x"4ac087c2",
   298 => x"5ac0d3c2",
   299 => x"87f1f126",
   300 => x"00000000",
   301 => x"00000000",
   302 => x"00000000",
   303 => x"00000000",
   304 => x"ff4a711e",
   305 => x"7249bfc8",
   306 => x"4f2648a1",
   307 => x"bfc8ff1e",
   308 => x"c0c0fe89",
   309 => x"a9c0c0c0",
   310 => x"c087c401",
   311 => x"c187c24a",
   312 => x"2648724a",
   313 => x"5b5e0e4f",
   314 => x"710e5d5c",
   315 => x"4cd4ff4b",
   316 => x"c04866d0",
   317 => x"ff49d678",
   318 => x"c387c5dc",
   319 => x"496c7cff",
   320 => x"7199ffc3",
   321 => x"f0c3494d",
   322 => x"a9e0c199",
   323 => x"c387cb05",
   324 => x"486c7cff",
   325 => x"66d098c3",
   326 => x"ffc37808",
   327 => x"494a6c7c",
   328 => x"ffc331c8",
   329 => x"714a6c7c",
   330 => x"c84972b2",
   331 => x"7cffc331",
   332 => x"b2714a6c",
   333 => x"31c84972",
   334 => x"6c7cffc3",
   335 => x"ffb2714a",
   336 => x"e0c048d0",
   337 => x"029b7378",
   338 => x"7b7287c2",
   339 => x"4d264875",
   340 => x"4b264c26",
   341 => x"261e4f26",
   342 => x"5b5e0e4f",
   343 => x"86f80e5c",
   344 => x"a6c81e76",
   345 => x"87fdfd49",
   346 => x"4b7086c4",
   347 => x"a8c4486e",
   348 => x"87f0c203",
   349 => x"f0c34a73",
   350 => x"aad0c19a",
   351 => x"c187c702",
   352 => x"c205aae0",
   353 => x"497387de",
   354 => x"c30299c8",
   355 => x"87c6ff87",
   356 => x"9cc34c73",
   357 => x"c105acc2",
   358 => x"66c487c2",
   359 => x"7131c949",
   360 => x"4a66c41e",
   361 => x"ecc292d4",
   362 => x"817249f1",
   363 => x"87d9d0fe",
   364 => x"d9ff49d8",
   365 => x"c0c887ca",
   366 => x"cedbc21e",
   367 => x"ddecfd49",
   368 => x"48d0ff87",
   369 => x"c278e0c0",
   370 => x"cc1ecedb",
   371 => x"92d44a66",
   372 => x"49f1ecc2",
   373 => x"cefe8172",
   374 => x"86cc87e1",
   375 => x"c105acc1",
   376 => x"66c487c2",
   377 => x"7131c949",
   378 => x"4a66c41e",
   379 => x"ecc292d4",
   380 => x"817249f1",
   381 => x"87d1cffe",
   382 => x"1ecedbc2",
   383 => x"d44a66c8",
   384 => x"f1ecc292",
   385 => x"fe817249",
   386 => x"d787e2cc",
   387 => x"efd7ff49",
   388 => x"1ec0c887",
   389 => x"49cedbc2",
   390 => x"87dbeafd",
   391 => x"d0ff86cc",
   392 => x"78e0c048",
   393 => x"e7fc8ef8",
   394 => x"5b5e0e87",
   395 => x"710e5d5c",
   396 => x"4cd4ff4a",
   397 => x"c34d66d0",
   398 => x"c506adb7",
   399 => x"c148c087",
   400 => x"1e7287e1",
   401 => x"93d44b75",
   402 => x"83f1ecc2",
   403 => x"c6fe4973",
   404 => x"83c887e7",
   405 => x"d0ff4b6b",
   406 => x"78e1c848",
   407 => x"48737cdd",
   408 => x"7098ffc3",
   409 => x"c849737c",
   410 => x"487129b7",
   411 => x"7098ffc3",
   412 => x"d049737c",
   413 => x"487129b7",
   414 => x"7098ffc3",
   415 => x"d848737c",
   416 => x"7c7028b7",
   417 => x"7c7c7cc0",
   418 => x"7c7c7c7c",
   419 => x"7c7c7c7c",
   420 => x"48d0ff7c",
   421 => x"7578e0c0",
   422 => x"ff49dc1e",
   423 => x"c887c6d6",
   424 => x"fa487386",
   425 => x"fa4887e8",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
