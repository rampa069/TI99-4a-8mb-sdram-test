
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"0c",x"18",x"0c",x"7c"),
     1 => (x"00",x"00",x"78",x"7c"),
     2 => (x"04",x"04",x"7c",x"7c"),
     3 => (x"00",x"00",x"78",x"7c"),
     4 => (x"44",x"44",x"7c",x"38"),
     5 => (x"00",x"00",x"38",x"7c"),
     6 => (x"24",x"24",x"fc",x"fc"),
     7 => (x"00",x"00",x"18",x"3c"),
     8 => (x"24",x"24",x"3c",x"18"),
     9 => (x"00",x"00",x"fc",x"fc"),
    10 => (x"04",x"04",x"7c",x"7c"),
    11 => (x"00",x"00",x"08",x"0c"),
    12 => (x"54",x"54",x"5c",x"48"),
    13 => (x"00",x"00",x"20",x"74"),
    14 => (x"44",x"7f",x"3f",x"04"),
    15 => (x"00",x"00",x"00",x"44"),
    16 => (x"40",x"40",x"7c",x"3c"),
    17 => (x"00",x"00",x"7c",x"7c"),
    18 => (x"60",x"60",x"3c",x"1c"),
    19 => (x"3c",x"00",x"1c",x"3c"),
    20 => (x"60",x"30",x"60",x"7c"),
    21 => (x"44",x"00",x"3c",x"7c"),
    22 => (x"38",x"10",x"38",x"6c"),
    23 => (x"00",x"00",x"44",x"6c"),
    24 => (x"60",x"e0",x"bc",x"1c"),
    25 => (x"00",x"00",x"1c",x"3c"),
    26 => (x"5c",x"74",x"64",x"44"),
    27 => (x"00",x"00",x"44",x"4c"),
    28 => (x"77",x"3e",x"08",x"08"),
    29 => (x"00",x"00",x"41",x"41"),
    30 => (x"7f",x"7f",x"00",x"00"),
    31 => (x"00",x"00",x"00",x"00"),
    32 => (x"3e",x"77",x"41",x"41"),
    33 => (x"02",x"00",x"08",x"08"),
    34 => (x"02",x"03",x"01",x"01"),
    35 => (x"7f",x"00",x"01",x"02"),
    36 => (x"7f",x"7f",x"7f",x"7f"),
    37 => (x"08",x"00",x"7f",x"7f"),
    38 => (x"3e",x"1c",x"1c",x"08"),
    39 => (x"7f",x"7f",x"7f",x"3e"),
    40 => (x"1c",x"3e",x"3e",x"7f"),
    41 => (x"00",x"08",x"08",x"1c"),
    42 => (x"7c",x"7c",x"18",x"10"),
    43 => (x"00",x"00",x"10",x"18"),
    44 => (x"7c",x"7c",x"30",x"10"),
    45 => (x"10",x"00",x"10",x"30"),
    46 => (x"78",x"60",x"60",x"30"),
    47 => (x"42",x"00",x"06",x"1e"),
    48 => (x"3c",x"18",x"3c",x"66"),
    49 => (x"78",x"00",x"42",x"66"),
    50 => (x"c6",x"c2",x"6a",x"38"),
    51 => (x"60",x"00",x"38",x"6c"),
    52 => (x"00",x"60",x"00",x"00"),
    53 => (x"0e",x"00",x"60",x"00"),
    54 => (x"5d",x"5c",x"5b",x"5e"),
    55 => (x"4c",x"71",x"1e",x"0e"),
    56 => (x"bf",x"e9",x"ec",x"c2"),
    57 => (x"c0",x"4b",x"c0",x"4d"),
    58 => (x"02",x"ab",x"74",x"1e"),
    59 => (x"a6",x"c4",x"87",x"c7"),
    60 => (x"c5",x"78",x"c0",x"48"),
    61 => (x"48",x"a6",x"c4",x"87"),
    62 => (x"66",x"c4",x"78",x"c1"),
    63 => (x"ee",x"49",x"73",x"1e"),
    64 => (x"86",x"c8",x"87",x"df"),
    65 => (x"ef",x"49",x"e0",x"c0"),
    66 => (x"a5",x"c4",x"87",x"ee"),
    67 => (x"f0",x"49",x"6a",x"4a"),
    68 => (x"c6",x"f1",x"87",x"f0"),
    69 => (x"c1",x"85",x"cb",x"87"),
    70 => (x"ab",x"b7",x"c8",x"83"),
    71 => (x"87",x"c7",x"ff",x"04"),
    72 => (x"26",x"4d",x"26",x"26"),
    73 => (x"26",x"4b",x"26",x"4c"),
    74 => (x"4a",x"71",x"1e",x"4f"),
    75 => (x"5a",x"ed",x"ec",x"c2"),
    76 => (x"48",x"ed",x"ec",x"c2"),
    77 => (x"fe",x"49",x"78",x"c7"),
    78 => (x"4f",x"26",x"87",x"dd"),
    79 => (x"71",x"1e",x"73",x"1e"),
    80 => (x"aa",x"b7",x"c0",x"4a"),
    81 => (x"c2",x"87",x"d3",x"03"),
    82 => (x"05",x"bf",x"f8",x"d2"),
    83 => (x"4b",x"c1",x"87",x"c4"),
    84 => (x"4b",x"c0",x"87",x"c2"),
    85 => (x"5b",x"fc",x"d2",x"c2"),
    86 => (x"d2",x"c2",x"87",x"c4"),
    87 => (x"d2",x"c2",x"5a",x"fc"),
    88 => (x"c1",x"4a",x"bf",x"f8"),
    89 => (x"a2",x"c0",x"c1",x"9a"),
    90 => (x"87",x"e8",x"ec",x"49"),
    91 => (x"d2",x"c2",x"48",x"fc"),
    92 => (x"fe",x"78",x"bf",x"f8"),
    93 => (x"71",x"1e",x"87",x"ef"),
    94 => (x"1e",x"66",x"c4",x"4a"),
    95 => (x"f9",x"ea",x"49",x"72"),
    96 => (x"4f",x"26",x"26",x"87"),
    97 => (x"48",x"d4",x"ff",x"1e"),
    98 => (x"ff",x"78",x"ff",x"c3"),
    99 => (x"e1",x"c0",x"48",x"d0"),
   100 => (x"48",x"d4",x"ff",x"78"),
   101 => (x"48",x"71",x"78",x"c1"),
   102 => (x"d4",x"ff",x"30",x"c4"),
   103 => (x"d0",x"ff",x"78",x"08"),
   104 => (x"78",x"e0",x"c0",x"48"),
   105 => (x"c2",x"1e",x"4f",x"26"),
   106 => (x"49",x"bf",x"f8",x"d2"),
   107 => (x"c2",x"87",x"f9",x"e6"),
   108 => (x"e8",x"48",x"e1",x"ec"),
   109 => (x"ec",x"c2",x"78",x"bf"),
   110 => (x"bf",x"ec",x"48",x"dd"),
   111 => (x"e1",x"ec",x"c2",x"78"),
   112 => (x"c3",x"49",x"4a",x"bf"),
   113 => (x"b7",x"c8",x"99",x"ff"),
   114 => (x"71",x"48",x"72",x"2a"),
   115 => (x"e9",x"ec",x"c2",x"b0"),
   116 => (x"0e",x"4f",x"26",x"58"),
   117 => (x"5d",x"5c",x"5b",x"5e"),
   118 => (x"ff",x"4b",x"71",x"0e"),
   119 => (x"ec",x"c2",x"87",x"c8"),
   120 => (x"50",x"c0",x"48",x"dc"),
   121 => (x"df",x"e6",x"49",x"73"),
   122 => (x"4c",x"49",x"70",x"87"),
   123 => (x"ee",x"cb",x"9c",x"c2"),
   124 => (x"87",x"cc",x"cb",x"49"),
   125 => (x"ec",x"c2",x"4d",x"70"),
   126 => (x"05",x"bf",x"97",x"dc"),
   127 => (x"d0",x"87",x"e2",x"c1"),
   128 => (x"ec",x"c2",x"49",x"66"),
   129 => (x"05",x"99",x"bf",x"e5"),
   130 => (x"66",x"d4",x"87",x"d6"),
   131 => (x"dd",x"ec",x"c2",x"49"),
   132 => (x"cb",x"05",x"99",x"bf"),
   133 => (x"e5",x"49",x"73",x"87"),
   134 => (x"98",x"70",x"87",x"ee"),
   135 => (x"87",x"c1",x"c1",x"02"),
   136 => (x"c1",x"fe",x"4c",x"c1"),
   137 => (x"ca",x"49",x"75",x"87"),
   138 => (x"98",x"70",x"87",x"e2"),
   139 => (x"c2",x"87",x"c6",x"02"),
   140 => (x"c1",x"48",x"dc",x"ec"),
   141 => (x"dc",x"ec",x"c2",x"50"),
   142 => (x"c0",x"05",x"bf",x"97"),
   143 => (x"ec",x"c2",x"87",x"e3"),
   144 => (x"d0",x"49",x"bf",x"e5"),
   145 => (x"ff",x"05",x"99",x"66"),
   146 => (x"ec",x"c2",x"87",x"d6"),
   147 => (x"d4",x"49",x"bf",x"dd"),
   148 => (x"ff",x"05",x"99",x"66"),
   149 => (x"49",x"73",x"87",x"ca"),
   150 => (x"70",x"87",x"ed",x"e4"),
   151 => (x"ff",x"fe",x"05",x"98"),
   152 => (x"fa",x"48",x"74",x"87"),
   153 => (x"5e",x"0e",x"87",x"fb"),
   154 => (x"0e",x"5d",x"5c",x"5b"),
   155 => (x"4d",x"c0",x"86",x"f8"),
   156 => (x"7e",x"bf",x"ec",x"4c"),
   157 => (x"c2",x"48",x"a6",x"c4"),
   158 => (x"78",x"bf",x"e9",x"ec"),
   159 => (x"1e",x"c0",x"1e",x"c1"),
   160 => (x"ce",x"fd",x"49",x"c7"),
   161 => (x"70",x"86",x"c8",x"87"),
   162 => (x"87",x"cd",x"02",x"98"),
   163 => (x"eb",x"fa",x"49",x"ff"),
   164 => (x"49",x"da",x"c1",x"87"),
   165 => (x"c1",x"87",x"f1",x"e3"),
   166 => (x"dc",x"ec",x"c2",x"4d"),
   167 => (x"cf",x"02",x"bf",x"97"),
   168 => (x"f0",x"d2",x"c2",x"87"),
   169 => (x"b9",x"c1",x"49",x"bf"),
   170 => (x"59",x"f4",x"d2",x"c2"),
   171 => (x"87",x"d4",x"fb",x"71"),
   172 => (x"bf",x"e1",x"ec",x"c2"),
   173 => (x"f8",x"d2",x"c2",x"4b"),
   174 => (x"e9",x"c0",x"05",x"bf"),
   175 => (x"49",x"fd",x"c3",x"87"),
   176 => (x"c3",x"87",x"c5",x"e3"),
   177 => (x"ff",x"e2",x"49",x"fa"),
   178 => (x"c3",x"49",x"73",x"87"),
   179 => (x"1e",x"71",x"99",x"ff"),
   180 => (x"e1",x"fa",x"49",x"c0"),
   181 => (x"c8",x"49",x"73",x"87"),
   182 => (x"1e",x"71",x"29",x"b7"),
   183 => (x"d5",x"fa",x"49",x"c1"),
   184 => (x"c5",x"86",x"c8",x"87"),
   185 => (x"ec",x"c2",x"87",x"f4"),
   186 => (x"9b",x"4b",x"bf",x"e5"),
   187 => (x"c2",x"87",x"dd",x"02"),
   188 => (x"49",x"bf",x"f4",x"d2"),
   189 => (x"70",x"87",x"d5",x"c7"),
   190 => (x"87",x"c4",x"05",x"98"),
   191 => (x"87",x"d2",x"4b",x"c0"),
   192 => (x"c6",x"49",x"e0",x"c2"),
   193 => (x"d2",x"c2",x"87",x"fa"),
   194 => (x"87",x"c6",x"58",x"f8"),
   195 => (x"48",x"f4",x"d2",x"c2"),
   196 => (x"49",x"73",x"78",x"c0"),
   197 => (x"cd",x"05",x"99",x"c2"),
   198 => (x"49",x"eb",x"c3",x"87"),
   199 => (x"70",x"87",x"e9",x"e1"),
   200 => (x"02",x"99",x"c2",x"49"),
   201 => (x"4c",x"fb",x"87",x"c2"),
   202 => (x"99",x"c1",x"49",x"73"),
   203 => (x"c3",x"87",x"cd",x"05"),
   204 => (x"d3",x"e1",x"49",x"f4"),
   205 => (x"c2",x"49",x"70",x"87"),
   206 => (x"87",x"c2",x"02",x"99"),
   207 => (x"49",x"73",x"4c",x"fa"),
   208 => (x"cd",x"05",x"99",x"c8"),
   209 => (x"49",x"f5",x"c3",x"87"),
   210 => (x"70",x"87",x"fd",x"e0"),
   211 => (x"02",x"99",x"c2",x"49"),
   212 => (x"ec",x"c2",x"87",x"d5"),
   213 => (x"ca",x"02",x"bf",x"ed"),
   214 => (x"88",x"c1",x"48",x"87"),
   215 => (x"58",x"f1",x"ec",x"c2"),
   216 => (x"ff",x"87",x"c2",x"c0"),
   217 => (x"73",x"4d",x"c1",x"4c"),
   218 => (x"05",x"99",x"c4",x"49"),
   219 => (x"f2",x"c3",x"87",x"cd"),
   220 => (x"87",x"d4",x"e0",x"49"),
   221 => (x"99",x"c2",x"49",x"70"),
   222 => (x"c2",x"87",x"dc",x"02"),
   223 => (x"7e",x"bf",x"ed",x"ec"),
   224 => (x"a8",x"b7",x"c7",x"48"),
   225 => (x"87",x"cb",x"c0",x"03"),
   226 => (x"80",x"c1",x"48",x"6e"),
   227 => (x"58",x"f1",x"ec",x"c2"),
   228 => (x"fe",x"87",x"c2",x"c0"),
   229 => (x"c3",x"4d",x"c1",x"4c"),
   230 => (x"df",x"ff",x"49",x"fd"),
   231 => (x"49",x"70",x"87",x"ea"),
   232 => (x"d5",x"02",x"99",x"c2"),
   233 => (x"ed",x"ec",x"c2",x"87"),
   234 => (x"c9",x"c0",x"02",x"bf"),
   235 => (x"ed",x"ec",x"c2",x"87"),
   236 => (x"c0",x"78",x"c0",x"48"),
   237 => (x"4c",x"fd",x"87",x"c2"),
   238 => (x"fa",x"c3",x"4d",x"c1"),
   239 => (x"c7",x"df",x"ff",x"49"),
   240 => (x"c2",x"49",x"70",x"87"),
   241 => (x"d9",x"c0",x"02",x"99"),
   242 => (x"ed",x"ec",x"c2",x"87"),
   243 => (x"b7",x"c7",x"48",x"bf"),
   244 => (x"c9",x"c0",x"03",x"a8"),
   245 => (x"ed",x"ec",x"c2",x"87"),
   246 => (x"c0",x"78",x"c7",x"48"),
   247 => (x"4c",x"fc",x"87",x"c2"),
   248 => (x"b7",x"c0",x"4d",x"c1"),
   249 => (x"d3",x"c0",x"03",x"ac"),
   250 => (x"48",x"66",x"c4",x"87"),
   251 => (x"70",x"80",x"d8",x"c1"),
   252 => (x"02",x"bf",x"6e",x"7e"),
   253 => (x"4b",x"87",x"c5",x"c0"),
   254 => (x"0f",x"73",x"49",x"74"),
   255 => (x"f0",x"c3",x"1e",x"c0"),
   256 => (x"49",x"da",x"c1",x"1e"),
   257 => (x"c8",x"87",x"cc",x"f7"),
   258 => (x"02",x"98",x"70",x"86"),
   259 => (x"c2",x"87",x"d8",x"c0"),
   260 => (x"7e",x"bf",x"ed",x"ec"),
   261 => (x"91",x"cb",x"49",x"6e"),
   262 => (x"71",x"4a",x"66",x"c4"),
   263 => (x"c0",x"02",x"6a",x"82"),
   264 => (x"6e",x"4b",x"87",x"c5"),
   265 => (x"75",x"0f",x"73",x"49"),
   266 => (x"c8",x"c0",x"02",x"9d"),
   267 => (x"ed",x"ec",x"c2",x"87"),
   268 => (x"e2",x"f2",x"49",x"bf"),
   269 => (x"fc",x"d2",x"c2",x"87"),
   270 => (x"dd",x"c0",x"02",x"bf"),
   271 => (x"cb",x"c2",x"49",x"87"),
   272 => (x"02",x"98",x"70",x"87"),
   273 => (x"c2",x"87",x"d3",x"c0"),
   274 => (x"49",x"bf",x"ed",x"ec"),
   275 => (x"c0",x"87",x"c8",x"f2"),
   276 => (x"87",x"e8",x"f3",x"49"),
   277 => (x"48",x"fc",x"d2",x"c2"),
   278 => (x"8e",x"f8",x"78",x"c0"),
   279 => (x"0e",x"87",x"c2",x"f3"),
   280 => (x"5d",x"5c",x"5b",x"5e"),
   281 => (x"4c",x"71",x"1e",x"0e"),
   282 => (x"bf",x"e9",x"ec",x"c2"),
   283 => (x"a1",x"cd",x"c1",x"49"),
   284 => (x"81",x"d1",x"c1",x"4d"),
   285 => (x"9c",x"74",x"7e",x"69"),
   286 => (x"c4",x"87",x"cf",x"02"),
   287 => (x"7b",x"74",x"4b",x"a5"),
   288 => (x"bf",x"e9",x"ec",x"c2"),
   289 => (x"87",x"e1",x"f2",x"49"),
   290 => (x"9c",x"74",x"7b",x"6e"),
   291 => (x"c0",x"87",x"c4",x"05"),
   292 => (x"c1",x"87",x"c2",x"4b"),
   293 => (x"f2",x"49",x"73",x"4b"),
   294 => (x"66",x"d4",x"87",x"e2"),
   295 => (x"49",x"87",x"c7",x"02"),
   296 => (x"4a",x"70",x"87",x"de"),
   297 => (x"4a",x"c0",x"87",x"c2"),
   298 => (x"5a",x"c0",x"d3",x"c2"),
   299 => (x"87",x"f1",x"f1",x"26"),
   300 => (x"00",x"00",x"00",x"00"),
   301 => (x"00",x"00",x"00",x"00"),
   302 => (x"00",x"00",x"00",x"00"),
   303 => (x"00",x"00",x"00",x"00"),
   304 => (x"ff",x"4a",x"71",x"1e"),
   305 => (x"72",x"49",x"bf",x"c8"),
   306 => (x"4f",x"26",x"48",x"a1"),
   307 => (x"bf",x"c8",x"ff",x"1e"),
   308 => (x"c0",x"c0",x"fe",x"89"),
   309 => (x"a9",x"c0",x"c0",x"c0"),
   310 => (x"c0",x"87",x"c4",x"01"),
   311 => (x"c1",x"87",x"c2",x"4a"),
   312 => (x"26",x"48",x"72",x"4a"),
   313 => (x"5b",x"5e",x"0e",x"4f"),
   314 => (x"71",x"0e",x"5d",x"5c"),
   315 => (x"4c",x"d4",x"ff",x"4b"),
   316 => (x"c0",x"48",x"66",x"d0"),
   317 => (x"ff",x"49",x"d6",x"78"),
   318 => (x"c3",x"87",x"c5",x"dc"),
   319 => (x"49",x"6c",x"7c",x"ff"),
   320 => (x"71",x"99",x"ff",x"c3"),
   321 => (x"f0",x"c3",x"49",x"4d"),
   322 => (x"a9",x"e0",x"c1",x"99"),
   323 => (x"c3",x"87",x"cb",x"05"),
   324 => (x"48",x"6c",x"7c",x"ff"),
   325 => (x"66",x"d0",x"98",x"c3"),
   326 => (x"ff",x"c3",x"78",x"08"),
   327 => (x"49",x"4a",x"6c",x"7c"),
   328 => (x"ff",x"c3",x"31",x"c8"),
   329 => (x"71",x"4a",x"6c",x"7c"),
   330 => (x"c8",x"49",x"72",x"b2"),
   331 => (x"7c",x"ff",x"c3",x"31"),
   332 => (x"b2",x"71",x"4a",x"6c"),
   333 => (x"31",x"c8",x"49",x"72"),
   334 => (x"6c",x"7c",x"ff",x"c3"),
   335 => (x"ff",x"b2",x"71",x"4a"),
   336 => (x"e0",x"c0",x"48",x"d0"),
   337 => (x"02",x"9b",x"73",x"78"),
   338 => (x"7b",x"72",x"87",x"c2"),
   339 => (x"4d",x"26",x"48",x"75"),
   340 => (x"4b",x"26",x"4c",x"26"),
   341 => (x"26",x"1e",x"4f",x"26"),
   342 => (x"5b",x"5e",x"0e",x"4f"),
   343 => (x"86",x"f8",x"0e",x"5c"),
   344 => (x"a6",x"c8",x"1e",x"76"),
   345 => (x"87",x"fd",x"fd",x"49"),
   346 => (x"4b",x"70",x"86",x"c4"),
   347 => (x"a8",x"c4",x"48",x"6e"),
   348 => (x"87",x"f0",x"c2",x"03"),
   349 => (x"f0",x"c3",x"4a",x"73"),
   350 => (x"aa",x"d0",x"c1",x"9a"),
   351 => (x"c1",x"87",x"c7",x"02"),
   352 => (x"c2",x"05",x"aa",x"e0"),
   353 => (x"49",x"73",x"87",x"de"),
   354 => (x"c3",x"02",x"99",x"c8"),
   355 => (x"87",x"c6",x"ff",x"87"),
   356 => (x"9c",x"c3",x"4c",x"73"),
   357 => (x"c1",x"05",x"ac",x"c2"),
   358 => (x"66",x"c4",x"87",x"c2"),
   359 => (x"71",x"31",x"c9",x"49"),
   360 => (x"4a",x"66",x"c4",x"1e"),
   361 => (x"ec",x"c2",x"92",x"d4"),
   362 => (x"81",x"72",x"49",x"f1"),
   363 => (x"87",x"d9",x"d0",x"fe"),
   364 => (x"d9",x"ff",x"49",x"d8"),
   365 => (x"c0",x"c8",x"87",x"ca"),
   366 => (x"ce",x"db",x"c2",x"1e"),
   367 => (x"dd",x"ec",x"fd",x"49"),
   368 => (x"48",x"d0",x"ff",x"87"),
   369 => (x"c2",x"78",x"e0",x"c0"),
   370 => (x"cc",x"1e",x"ce",x"db"),
   371 => (x"92",x"d4",x"4a",x"66"),
   372 => (x"49",x"f1",x"ec",x"c2"),
   373 => (x"ce",x"fe",x"81",x"72"),
   374 => (x"86",x"cc",x"87",x"e1"),
   375 => (x"c1",x"05",x"ac",x"c1"),
   376 => (x"66",x"c4",x"87",x"c2"),
   377 => (x"71",x"31",x"c9",x"49"),
   378 => (x"4a",x"66",x"c4",x"1e"),
   379 => (x"ec",x"c2",x"92",x"d4"),
   380 => (x"81",x"72",x"49",x"f1"),
   381 => (x"87",x"d1",x"cf",x"fe"),
   382 => (x"1e",x"ce",x"db",x"c2"),
   383 => (x"d4",x"4a",x"66",x"c8"),
   384 => (x"f1",x"ec",x"c2",x"92"),
   385 => (x"fe",x"81",x"72",x"49"),
   386 => (x"d7",x"87",x"e2",x"cc"),
   387 => (x"ef",x"d7",x"ff",x"49"),
   388 => (x"1e",x"c0",x"c8",x"87"),
   389 => (x"49",x"ce",x"db",x"c2"),
   390 => (x"87",x"db",x"ea",x"fd"),
   391 => (x"d0",x"ff",x"86",x"cc"),
   392 => (x"78",x"e0",x"c0",x"48"),
   393 => (x"e7",x"fc",x"8e",x"f8"),
   394 => (x"5b",x"5e",x"0e",x"87"),
   395 => (x"71",x"0e",x"5d",x"5c"),
   396 => (x"4c",x"d4",x"ff",x"4a"),
   397 => (x"c3",x"4d",x"66",x"d0"),
   398 => (x"c5",x"06",x"ad",x"b7"),
   399 => (x"c1",x"48",x"c0",x"87"),
   400 => (x"1e",x"72",x"87",x"e1"),
   401 => (x"93",x"d4",x"4b",x"75"),
   402 => (x"83",x"f1",x"ec",x"c2"),
   403 => (x"c6",x"fe",x"49",x"73"),
   404 => (x"83",x"c8",x"87",x"e7"),
   405 => (x"d0",x"ff",x"4b",x"6b"),
   406 => (x"78",x"e1",x"c8",x"48"),
   407 => (x"48",x"73",x"7c",x"dd"),
   408 => (x"70",x"98",x"ff",x"c3"),
   409 => (x"c8",x"49",x"73",x"7c"),
   410 => (x"48",x"71",x"29",x"b7"),
   411 => (x"70",x"98",x"ff",x"c3"),
   412 => (x"d0",x"49",x"73",x"7c"),
   413 => (x"48",x"71",x"29",x"b7"),
   414 => (x"70",x"98",x"ff",x"c3"),
   415 => (x"d8",x"48",x"73",x"7c"),
   416 => (x"7c",x"70",x"28",x"b7"),
   417 => (x"7c",x"7c",x"7c",x"c0"),
   418 => (x"7c",x"7c",x"7c",x"7c"),
   419 => (x"7c",x"7c",x"7c",x"7c"),
   420 => (x"48",x"d0",x"ff",x"7c"),
   421 => (x"75",x"78",x"e0",x"c0"),
   422 => (x"ff",x"49",x"dc",x"1e"),
   423 => (x"c8",x"87",x"c6",x"d6"),
   424 => (x"fa",x"48",x"73",x"86"),
   425 => (x"fa",x"48",x"87",x"e8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

