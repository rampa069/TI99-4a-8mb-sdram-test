library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8eec287",
    12 => x"86c0c84e",
    13 => x"49d8eec2",
    14 => x"48fcdac2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f4e2",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bffcda",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dac21e73",
   183 => x"78c148fc",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"c0dbc287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58c4dbc2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49c4dbc2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97c4db",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97cbdb",
   291 => x"c231d049",
   292 => x"bf97ccdb",
   293 => x"7232c84a",
   294 => x"cddbc2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dbc287e7",
   300 => x"49bf97cd",
   301 => x"99c631c1",
   302 => x"97cedbc2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97c9db",
   306 => x"9dcf4d4a",
   307 => x"97cadbc2",
   308 => x"9ac34abf",
   309 => x"dbc232ca",
   310 => x"4bbf97cb",
   311 => x"b27333c2",
   312 => x"97ccdbc2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e3c286f8",
   329 => x"78c048ea",
   330 => x"1ee2dbc2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"e2f2c07e",
   337 => x"dcc249bf",
   338 => x"c8714ad8",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfdef2",
   343 => x"4af4dcc2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e2c287fd",
   349 => x"c24dbfe8",
   350 => x"bf9fe0e3",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"e8e2c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"dbc287e3",
   359 => x"49751ee2",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfdef2",
   365 => x"4af4dcc2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148eae3",
   370 => x"c087da78",
   371 => x"49bfe2f2",
   372 => x"4ad8dcc2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"e0e3c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e3c287cd",
   381 => x"49bf97e1",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97e2dbc2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97eddbc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97eedb",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97efdbc2",
   400 => x"e3c248bf",
   401 => x"4c7058e6",
   402 => x"c288c148",
   403 => x"c258eae3",
   404 => x"bf97f0db",
   405 => x"c2817549",
   406 => x"bf97f1db",
   407 => x"7232c84a",
   408 => x"e7c27ea1",
   409 => x"786e48f7",
   410 => x"97f2dbc2",
   411 => x"a6c848bf",
   412 => x"eae3c258",
   413 => x"cfc202bf",
   414 => x"def2c087",
   415 => x"dcc249bf",
   416 => x"c8714af4",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbfe2e3",
   422 => x"5ccbe8c2",
   423 => x"97c7dcc2",
   424 => x"31c849bf",
   425 => x"97c6dcc2",
   426 => x"49a14abf",
   427 => x"97c8dcc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97c9dc",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"f7e7c291",
   434 => x"e7c281bf",
   435 => x"dcc259ff",
   436 => x"4abf97cf",
   437 => x"dcc232c8",
   438 => x"4bbf97ce",
   439 => x"dcc24aa2",
   440 => x"4bbf97d0",
   441 => x"a27333d0",
   442 => x"d1dcc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e8c24aa2",
   446 => x"8ac25ac3",
   447 => x"e8c29274",
   448 => x"a17248c3",
   449 => x"87c1c178",
   450 => x"97f4dbc2",
   451 => x"31c849bf",
   452 => x"97f3dbc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259cbe8",
   457 => x"bf97f9db",
   458 => x"c232c84a",
   459 => x"bf97f8db",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5ac7e8c2",
   463 => x"48ffe7c2",
   464 => x"e7c278c0",
   465 => x"a17248fb",
   466 => x"cbe8c278",
   467 => x"ffe7c248",
   468 => x"e8c278bf",
   469 => x"e8c248cf",
   470 => x"c278bfc3",
   471 => x"02bfeae3",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bfc7e8c2",
   476 => x"7030c448",
   477 => x"eee3c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfeae3",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e7c29dff",
   491 => x"c083bff7",
   492 => x"abbfdaf2",
   493 => x"c087d902",
   494 => x"c25bdef2",
   495 => x"731ee2db",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfeae3c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981e2db",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"e2dbc291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c1c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087eac2",
   521 => x"4949c11e",
   522 => x"c487d6ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4af2e3c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d4c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cfc102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfeae3",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"496e7ec0",
   556 => x"bf66c448",
   557 => x"0866c480",
   558 => x"cc7cc078",
   559 => x"66c449a4",
   560 => x"a4d079bf",
   561 => x"c179c049",
   562 => x"c087c248",
   563 => x"fa8ef848",
   564 => x"5e0e87ed",
   565 => x"0e5d5c5b",
   566 => x"029c4c71",
   567 => x"c887cbc1",
   568 => x"026949a4",
   569 => x"d087c3c1",
   570 => x"496c4a66",
   571 => x"7248a6d0",
   572 => x"b94d78a1",
   573 => x"bfe6e3c2",
   574 => x"72baff4a",
   575 => x"02997199",
   576 => x"c487e4c0",
   577 => x"496b4ba4",
   578 => x"7087fcf9",
   579 => x"e2e3c27b",
   580 => x"816c49bf",
   581 => x"b9757c71",
   582 => x"bfe6e3c2",
   583 => x"72baff4a",
   584 => x"05997199",
   585 => x"d087dcff",
   586 => x"d2f97c66",
   587 => x"1e731e87",
   588 => x"029b4b71",
   589 => x"a3c887c7",
   590 => x"c5056949",
   591 => x"c048c087",
   592 => x"e7c287f6",
   593 => x"c449bffb",
   594 => x"4a6a4aa3",
   595 => x"e3c28ac2",
   596 => x"7292bfe2",
   597 => x"e3c249a1",
   598 => x"6b4abfe6",
   599 => x"49a1729a",
   600 => x"59def2c0",
   601 => x"711e66c8",
   602 => x"c487e4ea",
   603 => x"05987086",
   604 => x"48c087c4",
   605 => x"48c187c2",
   606 => x"1e87c8f8",
   607 => x"4b711e73",
   608 => x"87c7029b",
   609 => x"6949a3c8",
   610 => x"c087c505",
   611 => x"87f6c048",
   612 => x"bffbe7c2",
   613 => x"4aa3c449",
   614 => x"8ac24a6a",
   615 => x"bfe2e3c2",
   616 => x"49a17292",
   617 => x"bfe6e3c2",
   618 => x"729a6b4a",
   619 => x"f2c049a1",
   620 => x"66c859de",
   621 => x"cfe6711e",
   622 => x"7086c487",
   623 => x"87c40598",
   624 => x"87c248c0",
   625 => x"faf648c1",
   626 => x"5b5e0e87",
   627 => x"1e0e5d5c",
   628 => x"66d44b71",
   629 => x"029b734d",
   630 => x"c887ccc1",
   631 => x"026949a3",
   632 => x"d087c4c1",
   633 => x"e3c24ca3",
   634 => x"ff49bfe6",
   635 => x"994a6cb9",
   636 => x"a966d47e",
   637 => x"c087cd06",
   638 => x"a3cc7c7b",
   639 => x"49a3c44a",
   640 => x"87ca796a",
   641 => x"c0f84972",
   642 => x"4d66d499",
   643 => x"49758d71",
   644 => x"1e7129c9",
   645 => x"f9fa4973",
   646 => x"e2dbc287",
   647 => x"fc49731e",
   648 => x"86c887cb",
   649 => x"267c66d4",
   650 => x"1e87d4f5",
   651 => x"4b711e73",
   652 => x"e4c0029b",
   653 => x"cfe8c287",
   654 => x"c24a735b",
   655 => x"e2e3c28a",
   656 => x"c29249bf",
   657 => x"48bffbe7",
   658 => x"e8c28072",
   659 => x"487158d3",
   660 => x"e3c230c4",
   661 => x"edc058f2",
   662 => x"cbe8c287",
   663 => x"ffe7c248",
   664 => x"e8c278bf",
   665 => x"e8c248cf",
   666 => x"c278bfc3",
   667 => x"02bfeae3",
   668 => x"e3c287c9",
   669 => x"c449bfe2",
   670 => x"c287c731",
   671 => x"49bfc7e8",
   672 => x"e3c231c4",
   673 => x"faf359f2",
   674 => x"5b5e0e87",
   675 => x"4a710e5c",
   676 => x"9a724bc0",
   677 => x"87e1c002",
   678 => x"9f49a2da",
   679 => x"e3c24b69",
   680 => x"cf02bfea",
   681 => x"49a2d487",
   682 => x"4c49699f",
   683 => x"9cffffc0",
   684 => x"87c234d0",
   685 => x"49744cc0",
   686 => x"fd4973b3",
   687 => x"c0f387ed",
   688 => x"5b5e0e87",
   689 => x"f40e5d5c",
   690 => x"c04a7186",
   691 => x"029a727e",
   692 => x"dbc287d8",
   693 => x"78c048de",
   694 => x"48d6dbc2",
   695 => x"bfcfe8c2",
   696 => x"dadbc278",
   697 => x"cbe8c248",
   698 => x"e3c278bf",
   699 => x"50c048ff",
   700 => x"bfeee3c2",
   701 => x"dedbc249",
   702 => x"aa714abf",
   703 => x"87c9c403",
   704 => x"99cf4972",
   705 => x"87e9c005",
   706 => x"48daf2c0",
   707 => x"bfd6dbc2",
   708 => x"e2dbc278",
   709 => x"d6dbc21e",
   710 => x"dbc249bf",
   711 => x"a1c148d6",
   712 => x"eae37178",
   713 => x"c086c487",
   714 => x"c248d6f2",
   715 => x"cc78e2db",
   716 => x"d6f2c087",
   717 => x"e0c048bf",
   718 => x"daf2c080",
   719 => x"dedbc258",
   720 => x"80c148bf",
   721 => x"58e2dbc2",
   722 => x"000c9627",
   723 => x"bf97bf00",
   724 => x"c2029d4d",
   725 => x"e5c387e3",
   726 => x"dcc202ad",
   727 => x"d6f2c087",
   728 => x"a3cb4bbf",
   729 => x"cf4c1149",
   730 => x"d2c105ac",
   731 => x"df497587",
   732 => x"cd89c199",
   733 => x"f2e3c291",
   734 => x"4aa3c181",
   735 => x"a3c35112",
   736 => x"c551124a",
   737 => x"51124aa3",
   738 => x"124aa3c7",
   739 => x"4aa3c951",
   740 => x"a3ce5112",
   741 => x"d051124a",
   742 => x"51124aa3",
   743 => x"124aa3d2",
   744 => x"4aa3d451",
   745 => x"a3d65112",
   746 => x"d851124a",
   747 => x"51124aa3",
   748 => x"124aa3dc",
   749 => x"4aa3de51",
   750 => x"7ec15112",
   751 => x"7487fac0",
   752 => x"0599c849",
   753 => x"7487ebc0",
   754 => x"0599d049",
   755 => x"66dc87d1",
   756 => x"87cbc002",
   757 => x"66dc4973",
   758 => x"0298700f",
   759 => x"6e87d3c0",
   760 => x"87c6c005",
   761 => x"48f2e3c2",
   762 => x"f2c050c0",
   763 => x"c248bfd6",
   764 => x"e3c287df",
   765 => x"50c048ff",
   766 => x"eee3c27e",
   767 => x"dbc249bf",
   768 => x"714abfde",
   769 => x"f7fb04aa",
   770 => x"cfe8c287",
   771 => x"c8c005bf",
   772 => x"eae3c287",
   773 => x"f6c102bf",
   774 => x"dadbc287",
   775 => x"e6ed49bf",
   776 => x"dedbc287",
   777 => x"48a6c458",
   778 => x"bfdadbc2",
   779 => x"eae3c278",
   780 => x"d8c002bf",
   781 => x"4966c487",
   782 => x"ffffffcf",
   783 => x"02a999f8",
   784 => x"c087c5c0",
   785 => x"87e1c04c",
   786 => x"dcc04cc1",
   787 => x"4966c487",
   788 => x"99f8ffcf",
   789 => x"c8c002a9",
   790 => x"48a6c887",
   791 => x"c5c078c0",
   792 => x"48a6c887",
   793 => x"66c878c1",
   794 => x"059c744c",
   795 => x"c487e0c0",
   796 => x"89c24966",
   797 => x"bfe2e3c2",
   798 => x"e7c2914a",
   799 => x"c24abffb",
   800 => x"7248d6db",
   801 => x"dbc278a1",
   802 => x"78c048de",
   803 => x"c087e1f9",
   804 => x"eb8ef448",
   805 => x"000087e9",
   806 => x"ffff0000",
   807 => x"0ca6ffff",
   808 => x"0caf0000",
   809 => x"41460000",
   810 => x"20323354",
   811 => x"46002020",
   812 => x"36315441",
   813 => x"00202020",
   814 => x"48d4ff1e",
   815 => x"6878ffc3",
   816 => x"1e4f2648",
   817 => x"c348d4ff",
   818 => x"d0ff78ff",
   819 => x"78e1c048",
   820 => x"d448d4ff",
   821 => x"d3e8c278",
   822 => x"bfd4ff48",
   823 => x"1e4f2650",
   824 => x"c048d0ff",
   825 => x"4f2678e0",
   826 => x"87ccff1e",
   827 => x"02994970",
   828 => x"fbc087c6",
   829 => x"87f105a9",
   830 => x"4f264871",
   831 => x"5c5b5e0e",
   832 => x"c04b710e",
   833 => x"87f0fe4c",
   834 => x"02994970",
   835 => x"c087f9c0",
   836 => x"c002a9ec",
   837 => x"fbc087f2",
   838 => x"ebc002a9",
   839 => x"b766cc87",
   840 => x"87c703ac",
   841 => x"c20266d0",
   842 => x"71537187",
   843 => x"87c20299",
   844 => x"c3fe84c1",
   845 => x"99497087",
   846 => x"c087cd02",
   847 => x"c702a9ec",
   848 => x"a9fbc087",
   849 => x"87d5ff05",
   850 => x"c30266d0",
   851 => x"7b97c087",
   852 => x"05a9ecc0",
   853 => x"4a7487c4",
   854 => x"4a7487c5",
   855 => x"728a0ac0",
   856 => x"2687c248",
   857 => x"264c264d",
   858 => x"1e4f264b",
   859 => x"7087c9fd",
   860 => x"aaf0c04a",
   861 => x"c087c904",
   862 => x"c301aaf9",
   863 => x"8af0c087",
   864 => x"04aac1c1",
   865 => x"dac187c9",
   866 => x"87c301aa",
   867 => x"728af7c0",
   868 => x"0e4f2648",
   869 => x"0e5c5b5e",
   870 => x"d4ff4a71",
   871 => x"c049724b",
   872 => x"4c7087e7",
   873 => x"87c2029c",
   874 => x"d0ff8cc1",
   875 => x"c178c548",
   876 => x"49747bd5",
   877 => x"e4c131c6",
   878 => x"4abf97d5",
   879 => x"70b07148",
   880 => x"48d0ff7b",
   881 => x"dcfe78c4",
   882 => x"5b5e0e87",
   883 => x"f80e5d5c",
   884 => x"c04c7186",
   885 => x"87ebfb7e",
   886 => x"f9c04bc0",
   887 => x"49bf97f6",
   888 => x"cf04a9c0",
   889 => x"87c0fc87",
   890 => x"f9c083c1",
   891 => x"49bf97f6",
   892 => x"87f106ab",
   893 => x"97f6f9c0",
   894 => x"87cf02bf",
   895 => x"7087f9fa",
   896 => x"c6029949",
   897 => x"a9ecc087",
   898 => x"c087f105",
   899 => x"87e8fa4b",
   900 => x"e3fa4d70",
   901 => x"58a6c887",
   902 => x"7087ddfa",
   903 => x"c883c14a",
   904 => x"699749a4",
   905 => x"c702ad49",
   906 => x"adffc087",
   907 => x"87e7c005",
   908 => x"9749a4c9",
   909 => x"66c44969",
   910 => x"87c702a9",
   911 => x"a8ffc048",
   912 => x"ca87d405",
   913 => x"699749a4",
   914 => x"c602aa49",
   915 => x"aaffc087",
   916 => x"c187c405",
   917 => x"c087d07e",
   918 => x"c602adec",
   919 => x"adfbc087",
   920 => x"c087c405",
   921 => x"6e7ec14b",
   922 => x"87e1fe02",
   923 => x"7387f0f9",
   924 => x"fb8ef848",
   925 => x"0e0087ed",
   926 => x"5d5c5b5e",
   927 => x"7186f80e",
   928 => x"4bd4ff4d",
   929 => x"e8c21e75",
   930 => x"ece549d8",
   931 => x"7086c487",
   932 => x"cac40298",
   933 => x"48a6c487",
   934 => x"bfd7e4c1",
   935 => x"fb497578",
   936 => x"d0ff87f1",
   937 => x"c178c548",
   938 => x"4ac07bd6",
   939 => x"1149a275",
   940 => x"cb82c17b",
   941 => x"f304aab7",
   942 => x"c34acc87",
   943 => x"82c17bff",
   944 => x"aab7e0c0",
   945 => x"ff87f404",
   946 => x"78c448d0",
   947 => x"c57bffc3",
   948 => x"7bd3c178",
   949 => x"78c47bc1",
   950 => x"b7c04866",
   951 => x"eec206a8",
   952 => x"e0e8c287",
   953 => x"66c44cbf",
   954 => x"c8887448",
   955 => x"9c7458a6",
   956 => x"87f7c102",
   957 => x"7ee2dbc2",
   958 => x"8c4dc0c8",
   959 => x"03acb7c0",
   960 => x"c0c887c6",
   961 => x"4cc04da4",
   962 => x"97d3e8c2",
   963 => x"99d049bf",
   964 => x"c087d002",
   965 => x"d8e8c21e",
   966 => x"87d1e849",
   967 => x"4a7086c4",
   968 => x"c287edc0",
   969 => x"c21ee2db",
   970 => x"e749d8e8",
   971 => x"86c487ff",
   972 => x"d0ff4a70",
   973 => x"78c5c848",
   974 => x"6e7bd4c1",
   975 => x"6e7bbf97",
   976 => x"7080c148",
   977 => x"058dc17e",
   978 => x"ff87f0ff",
   979 => x"78c448d0",
   980 => x"c5059a72",
   981 => x"c148c087",
   982 => x"1ec187c7",
   983 => x"49d8e8c2",
   984 => x"c487efe5",
   985 => x"059c7486",
   986 => x"c487c9fe",
   987 => x"b7c04866",
   988 => x"87d106a8",
   989 => x"48d8e8c2",
   990 => x"80d078c0",
   991 => x"80f478c0",
   992 => x"bfe4e8c2",
   993 => x"4866c478",
   994 => x"01a8b7c0",
   995 => x"ff87d2fd",
   996 => x"78c548d0",
   997 => x"c07bd3c1",
   998 => x"c178c47b",
   999 => x"c087c248",
  1000 => x"268ef848",
  1001 => x"264c264d",
  1002 => x"0e4f264b",
  1003 => x"5d5c5b5e",
  1004 => x"4b711e0e",
  1005 => x"ab4d4cc0",
  1006 => x"87e8c004",
  1007 => x"1ec9f7c0",
  1008 => x"c4029d75",
  1009 => x"c24ac087",
  1010 => x"724ac187",
  1011 => x"87f1eb49",
  1012 => x"7e7086c4",
  1013 => x"056e84c1",
  1014 => x"4c7387c2",
  1015 => x"ac7385c1",
  1016 => x"87d8ff06",
  1017 => x"fe26486e",
  1018 => x"5e0e87f9",
  1019 => x"710e5c5b",
  1020 => x"0266cc4b",
  1021 => x"c04c87d8",
  1022 => x"d8028cf0",
  1023 => x"c14a7487",
  1024 => x"87d1028a",
  1025 => x"87cd028a",
  1026 => x"87c9028a",
  1027 => x"497387d9",
  1028 => x"d287e4f9",
  1029 => x"c01e7487",
  1030 => x"d7d8c149",
  1031 => x"731e7487",
  1032 => x"cfd8c149",
  1033 => x"fd86c887",
  1034 => x"5e0e87fb",
  1035 => x"0e5d5c5b",
  1036 => x"494c711e",
  1037 => x"e9c291de",
  1038 => x"85714dc0",
  1039 => x"c1026d97",
  1040 => x"e8c287dc",
  1041 => x"7449bfec",
  1042 => x"defd7181",
  1043 => x"487e7087",
  1044 => x"f2c00298",
  1045 => x"f4e8c287",
  1046 => x"cb4a704b",
  1047 => x"c6c1ff49",
  1048 => x"cb4b7487",
  1049 => x"e9e4c193",
  1050 => x"c183c483",
  1051 => x"747be2c2",
  1052 => x"edc1c149",
  1053 => x"c17b7587",
  1054 => x"bf97d6e4",
  1055 => x"e8c21e49",
  1056 => x"e5fd49f4",
  1057 => x"7486c487",
  1058 => x"d5c1c149",
  1059 => x"c149c087",
  1060 => x"c287f4c2",
  1061 => x"c048d4e8",
  1062 => x"dd49c178",
  1063 => x"fc2687fb",
  1064 => x"6f4c87c1",
  1065 => x"6e696461",
  1066 => x"2e2e2e67",
  1067 => x"1e731e00",
  1068 => x"c2494a71",
  1069 => x"81bfece8",
  1070 => x"87effb71",
  1071 => x"029b4b70",
  1072 => x"e74987c4",
  1073 => x"e8c287c3",
  1074 => x"78c048ec",
  1075 => x"c8dd49c1",
  1076 => x"87d3fb87",
  1077 => x"c149c01e",
  1078 => x"2687ecc1",
  1079 => x"4a711e4f",
  1080 => x"c191cb49",
  1081 => x"c881e9e4",
  1082 => x"c2481181",
  1083 => x"c258d8e8",
  1084 => x"c048ece8",
  1085 => x"dc49c178",
  1086 => x"4f2687df",
  1087 => x"0299711e",
  1088 => x"e5c187d2",
  1089 => x"50c048fe",
  1090 => x"c3c180f7",
  1091 => x"e4c140dd",
  1092 => x"87ce78e2",
  1093 => x"48fae5c1",
  1094 => x"78dbe4c1",
  1095 => x"c3c180fc",
  1096 => x"4f2678d4",
  1097 => x"5c5b5e0e",
  1098 => x"86f40e5d",
  1099 => x"4de2dbc2",
  1100 => x"a6c44cc0",
  1101 => x"c278c048",
  1102 => x"48bfece8",
  1103 => x"c106a8c0",
  1104 => x"dbc287c0",
  1105 => x"029848e2",
  1106 => x"c087f7c0",
  1107 => x"c81ec9f7",
  1108 => x"87c70266",
  1109 => x"c048a6c4",
  1110 => x"c487c578",
  1111 => x"78c148a6",
  1112 => x"e54966c4",
  1113 => x"86c487db",
  1114 => x"84c14d70",
  1115 => x"c14866c4",
  1116 => x"58a6c880",
  1117 => x"bfece8c2",
  1118 => x"87c603ac",
  1119 => x"ff059d75",
  1120 => x"4cc087c9",
  1121 => x"c3029d75",
  1122 => x"f7c087dc",
  1123 => x"66c81ec9",
  1124 => x"cc87c702",
  1125 => x"78c048a6",
  1126 => x"a6cc87c5",
  1127 => x"cc78c148",
  1128 => x"dce44966",
  1129 => x"7086c487",
  1130 => x"0298487e",
  1131 => x"4987e4c2",
  1132 => x"699781cb",
  1133 => x"0299d049",
  1134 => x"7487d4c1",
  1135 => x"c191cb49",
  1136 => x"c181e9e4",
  1137 => x"c879edc2",
  1138 => x"51ffc381",
  1139 => x"91de4974",
  1140 => x"4dc0e9c2",
  1141 => x"c1c28571",
  1142 => x"a5c17d97",
  1143 => x"51e0c049",
  1144 => x"97f2e3c2",
  1145 => x"87d202bf",
  1146 => x"a5c284c1",
  1147 => x"f2e3c24b",
  1148 => x"fe49db4a",
  1149 => x"c187f0fa",
  1150 => x"a5cd87d9",
  1151 => x"c151c049",
  1152 => x"4ba5c284",
  1153 => x"49cb4a6e",
  1154 => x"87dbfafe",
  1155 => x"7487c4c1",
  1156 => x"c191cb49",
  1157 => x"c181e9e4",
  1158 => x"c279eac0",
  1159 => x"bf97f2e3",
  1160 => x"7487d802",
  1161 => x"c191de49",
  1162 => x"c0e9c284",
  1163 => x"c283714b",
  1164 => x"dd4af2e3",
  1165 => x"eef9fe49",
  1166 => x"7487d887",
  1167 => x"c293de4b",
  1168 => x"cb83c0e9",
  1169 => x"51c049a3",
  1170 => x"6e7384c1",
  1171 => x"fe49cb4a",
  1172 => x"c487d4f9",
  1173 => x"80c14866",
  1174 => x"c758a6c8",
  1175 => x"c5c003ac",
  1176 => x"fc056e87",
  1177 => x"487487e4",
  1178 => x"f6f48ef4",
  1179 => x"1e731e87",
  1180 => x"cb494b71",
  1181 => x"e9e4c191",
  1182 => x"4aa1c881",
  1183 => x"48d5e4c1",
  1184 => x"a1c95012",
  1185 => x"f6f9c04a",
  1186 => x"ca501248",
  1187 => x"d6e4c181",
  1188 => x"c1501148",
  1189 => x"bf97d6e4",
  1190 => x"49c01e49",
  1191 => x"c287cbf5",
  1192 => x"de48d4e8",
  1193 => x"d549c178",
  1194 => x"f32687ef",
  1195 => x"5e0e87f9",
  1196 => x"0e5d5c5b",
  1197 => x"4d7186f4",
  1198 => x"c191cb49",
  1199 => x"c881e9e4",
  1200 => x"a1ca4aa1",
  1201 => x"48a6c47e",
  1202 => x"bfdcecc2",
  1203 => x"bf976e78",
  1204 => x"4c66c44b",
  1205 => x"48122c73",
  1206 => x"7058a6cc",
  1207 => x"c984c19c",
  1208 => x"49699781",
  1209 => x"c204acb7",
  1210 => x"6e4cc087",
  1211 => x"c84abf97",
  1212 => x"31724966",
  1213 => x"66c4b9ff",
  1214 => x"72487499",
  1215 => x"484a7030",
  1216 => x"ecc2b071",
  1217 => x"e5c058e0",
  1218 => x"49c087d8",
  1219 => x"7587cad4",
  1220 => x"cdf7c049",
  1221 => x"f28ef487",
  1222 => x"731e87c9",
  1223 => x"494b711e",
  1224 => x"7387cbfe",
  1225 => x"87c6fe49",
  1226 => x"1e87fcf1",
  1227 => x"4b711e73",
  1228 => x"024aa3c6",
  1229 => x"8ac187db",
  1230 => x"8a87d602",
  1231 => x"87dac102",
  1232 => x"fcc0028a",
  1233 => x"c0028a87",
  1234 => x"028a87e1",
  1235 => x"dbc187cb",
  1236 => x"f649c787",
  1237 => x"dec187c7",
  1238 => x"ece8c287",
  1239 => x"cbc102bf",
  1240 => x"88c14887",
  1241 => x"58f0e8c2",
  1242 => x"c287c1c1",
  1243 => x"02bff0e8",
  1244 => x"c287f9c0",
  1245 => x"48bfece8",
  1246 => x"e8c280c1",
  1247 => x"ebc058f0",
  1248 => x"ece8c287",
  1249 => x"89c649bf",
  1250 => x"59f0e8c2",
  1251 => x"03a9b7c0",
  1252 => x"e8c287da",
  1253 => x"78c048ec",
  1254 => x"e8c287d2",
  1255 => x"cb02bff0",
  1256 => x"ece8c287",
  1257 => x"80c648bf",
  1258 => x"58f0e8c2",
  1259 => x"e8d149c0",
  1260 => x"c0497387",
  1261 => x"ef87ebf4",
  1262 => x"5e0e87ed",
  1263 => x"0e5d5c5b",
  1264 => x"dc86d4ff",
  1265 => x"a6c859a6",
  1266 => x"c478c048",
  1267 => x"66c0c180",
  1268 => x"c180c478",
  1269 => x"c180c478",
  1270 => x"f0e8c278",
  1271 => x"c278c148",
  1272 => x"48bfd4e8",
  1273 => x"c905a8de",
  1274 => x"87f8f487",
  1275 => x"cf58a6cc",
  1276 => x"cee387e6",
  1277 => x"87f0e387",
  1278 => x"7087fde2",
  1279 => x"acfbc04c",
  1280 => x"87fbc102",
  1281 => x"c10566d8",
  1282 => x"fcc087ed",
  1283 => x"82c44a66",
  1284 => x"1e727e6a",
  1285 => x"48cde0c1",
  1286 => x"c84966c4",
  1287 => x"41204aa1",
  1288 => x"f905aa71",
  1289 => x"26511087",
  1290 => x"66fcc04a",
  1291 => x"edc9c148",
  1292 => x"c7496a78",
  1293 => x"c0517481",
  1294 => x"c84966fc",
  1295 => x"c051c181",
  1296 => x"c94966fc",
  1297 => x"c051c081",
  1298 => x"ca4966fc",
  1299 => x"c151c081",
  1300 => x"6a1ed81e",
  1301 => x"e281c849",
  1302 => x"86c887e2",
  1303 => x"4866c0c1",
  1304 => x"c701a8c0",
  1305 => x"48a6c887",
  1306 => x"87ce78c1",
  1307 => x"4866c0c1",
  1308 => x"a6d088c1",
  1309 => x"e187c358",
  1310 => x"a6d087ee",
  1311 => x"7478c248",
  1312 => x"cfcd029c",
  1313 => x"4866c887",
  1314 => x"a866c4c1",
  1315 => x"87c4cd03",
  1316 => x"c048a6dc",
  1317 => x"c080e878",
  1318 => x"87dce078",
  1319 => x"d0c14c70",
  1320 => x"d7c205ac",
  1321 => x"7e66c487",
  1322 => x"c887c0e3",
  1323 => x"c7e058a6",
  1324 => x"c04c7087",
  1325 => x"c105acec",
  1326 => x"66c887ed",
  1327 => x"c091cb49",
  1328 => x"c48166fc",
  1329 => x"4d6a4aa1",
  1330 => x"c44aa1c8",
  1331 => x"c3c15266",
  1332 => x"dfff79dd",
  1333 => x"4c7087e2",
  1334 => x"87d9029c",
  1335 => x"02acfbc0",
  1336 => x"557487d3",
  1337 => x"87d0dfff",
  1338 => x"029c4c70",
  1339 => x"fbc087c7",
  1340 => x"edff05ac",
  1341 => x"55e0c087",
  1342 => x"c055c1c2",
  1343 => x"66d87d97",
  1344 => x"05a86e48",
  1345 => x"66c887db",
  1346 => x"a866cc48",
  1347 => x"c887ca04",
  1348 => x"80c14866",
  1349 => x"c858a6cc",
  1350 => x"4866cc87",
  1351 => x"a6d088c1",
  1352 => x"d3deff58",
  1353 => x"c14c7087",
  1354 => x"c805acd0",
  1355 => x"4866d487",
  1356 => x"a6d880c1",
  1357 => x"acd0c158",
  1358 => x"87e9fd02",
  1359 => x"d84866c4",
  1360 => x"c905a866",
  1361 => x"e0c087e0",
  1362 => x"78c048a6",
  1363 => x"fbc04874",
  1364 => x"487e7088",
  1365 => x"e2c90298",
  1366 => x"88cb4887",
  1367 => x"98487e70",
  1368 => x"87cdc102",
  1369 => x"7088c948",
  1370 => x"0298487e",
  1371 => x"4887fec3",
  1372 => x"7e7088c4",
  1373 => x"ce029848",
  1374 => x"88c14887",
  1375 => x"98487e70",
  1376 => x"87e9c302",
  1377 => x"dc87d6c8",
  1378 => x"f0c048a6",
  1379 => x"e7dcff78",
  1380 => x"c04c7087",
  1381 => x"c002acec",
  1382 => x"e0c087c4",
  1383 => x"ecc05ca6",
  1384 => x"87cd02ac",
  1385 => x"87d0dcff",
  1386 => x"ecc04c70",
  1387 => x"f3ff05ac",
  1388 => x"acecc087",
  1389 => x"87c4c002",
  1390 => x"87fcdbff",
  1391 => x"1eca1ec0",
  1392 => x"cb4966d0",
  1393 => x"66c4c191",
  1394 => x"cc807148",
  1395 => x"66c858a6",
  1396 => x"d080c448",
  1397 => x"66cc58a6",
  1398 => x"dcff49bf",
  1399 => x"1ec187de",
  1400 => x"66d41ede",
  1401 => x"dcff49bf",
  1402 => x"86d087d2",
  1403 => x"c0484970",
  1404 => x"e8c08808",
  1405 => x"a8c058a6",
  1406 => x"87eec006",
  1407 => x"4866e4c0",
  1408 => x"c003a8dd",
  1409 => x"66c487e4",
  1410 => x"e4c049bf",
  1411 => x"e0c08166",
  1412 => x"66e4c051",
  1413 => x"c481c149",
  1414 => x"c281bf66",
  1415 => x"e4c051c1",
  1416 => x"81c24966",
  1417 => x"81bf66c4",
  1418 => x"486e51c0",
  1419 => x"78edc9c1",
  1420 => x"81c8496e",
  1421 => x"6e5166d0",
  1422 => x"d481c949",
  1423 => x"496e5166",
  1424 => x"66dc81ca",
  1425 => x"4866d051",
  1426 => x"a6d480c1",
  1427 => x"4866c858",
  1428 => x"04a866cc",
  1429 => x"c887cbc0",
  1430 => x"80c14866",
  1431 => x"c558a6cc",
  1432 => x"66cc87d9",
  1433 => x"d088c148",
  1434 => x"cec558a6",
  1435 => x"fadbff87",
  1436 => x"a6e8c087",
  1437 => x"f2dbff58",
  1438 => x"a6e0c087",
  1439 => x"a8ecc058",
  1440 => x"87cac005",
  1441 => x"c048a6dc",
  1442 => x"c07866e4",
  1443 => x"d8ff87c4",
  1444 => x"66c887e6",
  1445 => x"c091cb49",
  1446 => x"714866fc",
  1447 => x"4a7e7080",
  1448 => x"496e82c8",
  1449 => x"e4c081ca",
  1450 => x"66dc5166",
  1451 => x"c081c149",
  1452 => x"c18966e4",
  1453 => x"70307148",
  1454 => x"7189c149",
  1455 => x"ecc27a97",
  1456 => x"c049bfdc",
  1457 => x"972966e4",
  1458 => x"71484a6a",
  1459 => x"a6ecc098",
  1460 => x"c4496e58",
  1461 => x"d84d6981",
  1462 => x"66c44866",
  1463 => x"c8c002a8",
  1464 => x"48a6c487",
  1465 => x"c5c078c0",
  1466 => x"48a6c487",
  1467 => x"66c478c1",
  1468 => x"1ee0c01e",
  1469 => x"d8ff4975",
  1470 => x"86c887c2",
  1471 => x"b7c04c70",
  1472 => x"d4c106ac",
  1473 => x"c0857487",
  1474 => x"897449e0",
  1475 => x"e0c14b75",
  1476 => x"fe714ad6",
  1477 => x"c287d0e6",
  1478 => x"66e0c085",
  1479 => x"c080c148",
  1480 => x"c058a6e4",
  1481 => x"c14966e8",
  1482 => x"02a97081",
  1483 => x"c487c8c0",
  1484 => x"78c048a6",
  1485 => x"c487c5c0",
  1486 => x"78c148a6",
  1487 => x"c21e66c4",
  1488 => x"e0c049a4",
  1489 => x"70887148",
  1490 => x"49751e49",
  1491 => x"87ecd6ff",
  1492 => x"b7c086c8",
  1493 => x"c0ff01a8",
  1494 => x"66e0c087",
  1495 => x"87d1c002",
  1496 => x"81c9496e",
  1497 => x"5166e0c0",
  1498 => x"cac1486e",
  1499 => x"ccc078ee",
  1500 => x"c9496e87",
  1501 => x"6e51c281",
  1502 => x"daccc148",
  1503 => x"4866c878",
  1504 => x"04a866cc",
  1505 => x"c887cbc0",
  1506 => x"80c14866",
  1507 => x"c058a6cc",
  1508 => x"66cc87e9",
  1509 => x"d088c148",
  1510 => x"dec058a6",
  1511 => x"c7d5ff87",
  1512 => x"c04c7087",
  1513 => x"c6c187d5",
  1514 => x"c8c005ac",
  1515 => x"4866d087",
  1516 => x"a6d480c1",
  1517 => x"efd4ff58",
  1518 => x"d44c7087",
  1519 => x"80c14866",
  1520 => x"7458a6d8",
  1521 => x"cbc0029c",
  1522 => x"4866c887",
  1523 => x"a866c4c1",
  1524 => x"87fcf204",
  1525 => x"87c7d4ff",
  1526 => x"c74866c8",
  1527 => x"e5c003a8",
  1528 => x"f0e8c287",
  1529 => x"c878c048",
  1530 => x"91cb4966",
  1531 => x"8166fcc0",
  1532 => x"6a4aa1c4",
  1533 => x"7952c04a",
  1534 => x"c14866c8",
  1535 => x"58a6cc80",
  1536 => x"ff04a8c7",
  1537 => x"d4ff87db",
  1538 => x"d6deff8e",
  1539 => x"616f4c87",
  1540 => x"2e2a2064",
  1541 => x"203a0020",
  1542 => x"1e731e00",
  1543 => x"029b4b71",
  1544 => x"e8c287c6",
  1545 => x"78c048ec",
  1546 => x"e8c21ec7",
  1547 => x"c11ebfec",
  1548 => x"c21ee9e4",
  1549 => x"49bfd4e8",
  1550 => x"cc87ffed",
  1551 => x"d4e8c286",
  1552 => x"f7e249bf",
  1553 => x"029b7387",
  1554 => x"e4c187c8",
  1555 => x"e3c049e9",
  1556 => x"ddff87e2",
  1557 => x"731e87d1",
  1558 => x"c14bc01e",
  1559 => x"c048d5e4",
  1560 => x"cce6c150",
  1561 => x"d8ff49bf",
  1562 => x"987087cd",
  1563 => x"c187c405",
  1564 => x"734bf9e1",
  1565 => x"eedcff48",
  1566 => x"4d4f5287",
  1567 => x"616f6c20",
  1568 => x"676e6964",
  1569 => x"69616620",
  1570 => x"0064656c",
  1571 => x"87e3c71e",
  1572 => x"c4fe49c1",
  1573 => x"fee8fe87",
  1574 => x"02987087",
  1575 => x"f1fe87cd",
  1576 => x"987087f8",
  1577 => x"c187c402",
  1578 => x"c087c24a",
  1579 => x"059a724a",
  1580 => x"1ec087ce",
  1581 => x"49dce3c1",
  1582 => x"87eeeec0",
  1583 => x"87fe86c4",
  1584 => x"e3c11ec0",
  1585 => x"eec049e7",
  1586 => x"1ec087e0",
  1587 => x"7087c7fe",
  1588 => x"d5eec049",
  1589 => x"87dac387",
  1590 => x"4f268ef8",
  1591 => x"66204453",
  1592 => x"656c6961",
  1593 => x"42002e64",
  1594 => x"69746f6f",
  1595 => x"2e2e676e",
  1596 => x"c01e002e",
  1597 => x"c087fae5",
  1598 => x"f687e9f1",
  1599 => x"1e4f2687",
  1600 => x"48ece8c2",
  1601 => x"e8c278c0",
  1602 => x"78c048d4",
  1603 => x"e187fdfd",
  1604 => x"2648c087",
  1605 => x"0100004f",
  1606 => x"80000000",
  1607 => x"69784520",
  1608 => x"20800074",
  1609 => x"6b636142",
  1610 => x"00102a00",
  1611 => x"002a4000",
  1612 => x"00000000",
  1613 => x"0000102a",
  1614 => x"00002a5e",
  1615 => x"2a000000",
  1616 => x"7c000010",
  1617 => x"0000002a",
  1618 => x"102a0000",
  1619 => x"2a9a0000",
  1620 => x"00000000",
  1621 => x"00102a00",
  1622 => x"002ab800",
  1623 => x"00000000",
  1624 => x"0000102a",
  1625 => x"00002ad6",
  1626 => x"2a000000",
  1627 => x"f4000010",
  1628 => x"0000002a",
  1629 => x"10dd0000",
  1630 => x"00000000",
  1631 => x"00000000",
  1632 => x"00132b00",
  1633 => x"00000000",
  1634 => x"00000000",
  1635 => x"00001990",
  1636 => x"39394954",
  1637 => x"20204134",
  1638 => x"004d4f52",
  1639 => x"48f0fe1e",
  1640 => x"09cd78c0",
  1641 => x"4f260979",
  1642 => x"f0fe1e1e",
  1643 => x"26487ebf",
  1644 => x"fe1e4f26",
  1645 => x"78c148f0",
  1646 => x"fe1e4f26",
  1647 => x"78c048f0",
  1648 => x"711e4f26",
  1649 => x"5252c04a",
  1650 => x"5e0e4f26",
  1651 => x"0e5d5c5b",
  1652 => x"4d7186f4",
  1653 => x"c17e6d97",
  1654 => x"6c974ca5",
  1655 => x"58a6c848",
  1656 => x"66c4486e",
  1657 => x"87c505a8",
  1658 => x"e6c048ff",
  1659 => x"87caff87",
  1660 => x"9749a5c2",
  1661 => x"a3714b6c",
  1662 => x"4b6b974b",
  1663 => x"6e7e6c97",
  1664 => x"c880c148",
  1665 => x"98c758a6",
  1666 => x"7058a6cc",
  1667 => x"e1fe7c97",
  1668 => x"f4487387",
  1669 => x"264d268e",
  1670 => x"264b264c",
  1671 => x"5b5e0e4f",
  1672 => x"86f40e5c",
  1673 => x"66d84c71",
  1674 => x"9affc34a",
  1675 => x"974ba4c2",
  1676 => x"a173496c",
  1677 => x"97517249",
  1678 => x"486e7e6c",
  1679 => x"a6c880c1",
  1680 => x"cc98c758",
  1681 => x"547058a6",
  1682 => x"caff8ef4",
  1683 => x"fd1e1e87",
  1684 => x"bfe087e8",
  1685 => x"e0c0494a",
  1686 => x"cb0299c0",
  1687 => x"c21e7287",
  1688 => x"fe49d2ec",
  1689 => x"86c487f7",
  1690 => x"7087fdfc",
  1691 => x"87c2fd7e",
  1692 => x"1e4f2626",
  1693 => x"49d2ecc2",
  1694 => x"c187c7fd",
  1695 => x"fc49cde9",
  1696 => x"f7c387da",
  1697 => x"0e4f2687",
  1698 => x"5d5c5b5e",
  1699 => x"c24d710e",
  1700 => x"fc49d2ec",
  1701 => x"4b7087f4",
  1702 => x"04abb7c0",
  1703 => x"c387c2c3",
  1704 => x"c905abf0",
  1705 => x"ebedc187",
  1706 => x"c278c148",
  1707 => x"e0c387e3",
  1708 => x"87c905ab",
  1709 => x"48efedc1",
  1710 => x"d4c278c1",
  1711 => x"efedc187",
  1712 => x"87c602bf",
  1713 => x"4ca3c0c2",
  1714 => x"4c7387c2",
  1715 => x"bfebedc1",
  1716 => x"87e0c002",
  1717 => x"b7c44974",
  1718 => x"efc19129",
  1719 => x"4a7481cb",
  1720 => x"92c29acf",
  1721 => x"307248c1",
  1722 => x"baff4a70",
  1723 => x"98694872",
  1724 => x"87db7970",
  1725 => x"b7c44974",
  1726 => x"efc19129",
  1727 => x"4a7481cb",
  1728 => x"92c29acf",
  1729 => x"307248c3",
  1730 => x"69484a70",
  1731 => x"757970b0",
  1732 => x"f0c0059d",
  1733 => x"48d0ff87",
  1734 => x"ff78e1c8",
  1735 => x"78c548d4",
  1736 => x"bfefedc1",
  1737 => x"c387c302",
  1738 => x"edc178e0",
  1739 => x"c602bfeb",
  1740 => x"48d4ff87",
  1741 => x"ff78f0c3",
  1742 => x"0b7b0bd4",
  1743 => x"c848d0ff",
  1744 => x"e0c078e1",
  1745 => x"efedc178",
  1746 => x"c178c048",
  1747 => x"c048ebed",
  1748 => x"d2ecc278",
  1749 => x"87f2f949",
  1750 => x"b7c04b70",
  1751 => x"fefc03ab",
  1752 => x"2648c087",
  1753 => x"264c264d",
  1754 => x"004f264b",
  1755 => x"00000000",
  1756 => x"1e000000",
  1757 => x"fc494a71",
  1758 => x"4f2687cd",
  1759 => x"724ac01e",
  1760 => x"c191c449",
  1761 => x"c081cbef",
  1762 => x"d082c179",
  1763 => x"ee04aab7",
  1764 => x"0e4f2687",
  1765 => x"5d5c5b5e",
  1766 => x"f84d710e",
  1767 => x"4a7587dc",
  1768 => x"922ab7c4",
  1769 => x"82cbefc1",
  1770 => x"9ccf4c75",
  1771 => x"496a94c2",
  1772 => x"c32b744b",
  1773 => x"7448c29b",
  1774 => x"ff4c7030",
  1775 => x"714874bc",
  1776 => x"f77a7098",
  1777 => x"487387ec",
  1778 => x"0087d8fe",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"1e000000",
  1795 => x"c848d0ff",
  1796 => x"487178e1",
  1797 => x"7808d4ff",
  1798 => x"ff1e4f26",
  1799 => x"e1c848d0",
  1800 => x"ff487178",
  1801 => x"c47808d4",
  1802 => x"d4ff4866",
  1803 => x"4f267808",
  1804 => x"c44a711e",
  1805 => x"721e4966",
  1806 => x"87deff49",
  1807 => x"c048d0ff",
  1808 => x"262678e0",
  1809 => x"1e731e4f",
  1810 => x"66c84b71",
  1811 => x"4a731e49",
  1812 => x"49a2e0c1",
  1813 => x"2687d9ff",
  1814 => x"4d2687c4",
  1815 => x"4b264c26",
  1816 => x"ff1e4f26",
  1817 => x"ffc34ad4",
  1818 => x"48d0ff7a",
  1819 => x"de78e1c0",
  1820 => x"dcecc27a",
  1821 => x"48497abf",
  1822 => x"7a7028c8",
  1823 => x"28d04871",
  1824 => x"48717a70",
  1825 => x"7a7028d8",
  1826 => x"c048d0ff",
  1827 => x"4f2678e0",
  1828 => x"48d0ff1e",
  1829 => x"7178c9c8",
  1830 => x"08d4ff48",
  1831 => x"1e4f2678",
  1832 => x"eb494a71",
  1833 => x"48d0ff87",
  1834 => x"4f2678c8",
  1835 => x"711e731e",
  1836 => x"ececc24b",
  1837 => x"87c302bf",
  1838 => x"ff87ebc2",
  1839 => x"c9c848d0",
  1840 => x"c0487378",
  1841 => x"d4ffb0e0",
  1842 => x"ecc27808",
  1843 => x"78c048e0",
  1844 => x"c50266c8",
  1845 => x"49ffc387",
  1846 => x"49c087c2",
  1847 => x"59e8ecc2",
  1848 => x"c60266cc",
  1849 => x"d5d5c587",
  1850 => x"cf87c44a",
  1851 => x"c24affff",
  1852 => x"c25aecec",
  1853 => x"c148ecec",
  1854 => x"2687c478",
  1855 => x"264c264d",
  1856 => x"0e4f264b",
  1857 => x"5d5c5b5e",
  1858 => x"c24a710e",
  1859 => x"4cbfe8ec",
  1860 => x"cb029a72",
  1861 => x"91c84987",
  1862 => x"4be2f2c1",
  1863 => x"87c48371",
  1864 => x"4be2f6c1",
  1865 => x"49134dc0",
  1866 => x"ecc29974",
  1867 => x"7148bfe4",
  1868 => x"08d4ffb8",
  1869 => x"2cb7c178",
  1870 => x"adb7c885",
  1871 => x"c287e704",
  1872 => x"48bfe0ec",
  1873 => x"ecc280c8",
  1874 => x"eefe58e4",
  1875 => x"1e731e87",
  1876 => x"4a134b71",
  1877 => x"87cb029a",
  1878 => x"e6fe4972",
  1879 => x"9a4a1387",
  1880 => x"fe87f505",
  1881 => x"c21e87d9",
  1882 => x"49bfe0ec",
  1883 => x"48e0ecc2",
  1884 => x"c478a1c1",
  1885 => x"03a9b7c0",
  1886 => x"d4ff87db",
  1887 => x"e4ecc248",
  1888 => x"ecc278bf",
  1889 => x"c249bfe0",
  1890 => x"c148e0ec",
  1891 => x"c0c478a1",
  1892 => x"e504a9b7",
  1893 => x"48d0ff87",
  1894 => x"ecc278c8",
  1895 => x"78c048ec",
  1896 => x"00004f26",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"005f5f00",
  1900 => x"03000000",
  1901 => x"03030003",
  1902 => x"7f140000",
  1903 => x"7f7f147f",
  1904 => x"24000014",
  1905 => x"3a6b6b2e",
  1906 => x"6a4c0012",
  1907 => x"566c1836",
  1908 => x"7e300032",
  1909 => x"3a77594f",
  1910 => x"00004068",
  1911 => x"00030704",
  1912 => x"00000000",
  1913 => x"41633e1c",
  1914 => x"00000000",
  1915 => x"1c3e6341",
  1916 => x"2a080000",
  1917 => x"3e1c1c3e",
  1918 => x"0800082a",
  1919 => x"083e3e08",
  1920 => x"00000008",
  1921 => x"0060e080",
  1922 => x"08000000",
  1923 => x"08080808",
  1924 => x"00000008",
  1925 => x"00606000",
  1926 => x"60400000",
  1927 => x"060c1830",
  1928 => x"3e000103",
  1929 => x"7f4d597f",
  1930 => x"0400003e",
  1931 => x"007f7f06",
  1932 => x"42000000",
  1933 => x"4f597163",
  1934 => x"22000046",
  1935 => x"7f494963",
  1936 => x"1c180036",
  1937 => x"7f7f1316",
  1938 => x"27000010",
  1939 => x"7d454567",
  1940 => x"3c000039",
  1941 => x"79494b7e",
  1942 => x"01000030",
  1943 => x"0f797101",
  1944 => x"36000007",
  1945 => x"7f49497f",
  1946 => x"06000036",
  1947 => x"3f69494f",
  1948 => x"0000001e",
  1949 => x"00666600",
  1950 => x"00000000",
  1951 => x"0066e680",
  1952 => x"08000000",
  1953 => x"22141408",
  1954 => x"14000022",
  1955 => x"14141414",
  1956 => x"22000014",
  1957 => x"08141422",
  1958 => x"02000008",
  1959 => x"0f595103",
  1960 => x"7f3e0006",
  1961 => x"1f555d41",
  1962 => x"7e00001e",
  1963 => x"7f09097f",
  1964 => x"7f00007e",
  1965 => x"7f49497f",
  1966 => x"1c000036",
  1967 => x"4141633e",
  1968 => x"7f000041",
  1969 => x"3e63417f",
  1970 => x"7f00001c",
  1971 => x"4149497f",
  1972 => x"7f000041",
  1973 => x"0109097f",
  1974 => x"3e000001",
  1975 => x"7b49417f",
  1976 => x"7f00007a",
  1977 => x"7f08087f",
  1978 => x"0000007f",
  1979 => x"417f7f41",
  1980 => x"20000000",
  1981 => x"7f404060",
  1982 => x"7f7f003f",
  1983 => x"63361c08",
  1984 => x"7f000041",
  1985 => x"4040407f",
  1986 => x"7f7f0040",
  1987 => x"7f060c06",
  1988 => x"7f7f007f",
  1989 => x"7f180c06",
  1990 => x"3e00007f",
  1991 => x"7f41417f",
  1992 => x"7f00003e",
  1993 => x"0f09097f",
  1994 => x"7f3e0006",
  1995 => x"7e7f6141",
  1996 => x"7f000040",
  1997 => x"7f19097f",
  1998 => x"26000066",
  1999 => x"7b594d6f",
  2000 => x"01000032",
  2001 => x"017f7f01",
  2002 => x"3f000001",
  2003 => x"7f40407f",
  2004 => x"0f00003f",
  2005 => x"3f70703f",
  2006 => x"7f7f000f",
  2007 => x"7f301830",
  2008 => x"6341007f",
  2009 => x"361c1c36",
  2010 => x"03014163",
  2011 => x"067c7c06",
  2012 => x"71610103",
  2013 => x"43474d59",
  2014 => x"00000041",
  2015 => x"41417f7f",
  2016 => x"03010000",
  2017 => x"30180c06",
  2018 => x"00004060",
  2019 => x"7f7f4141",
  2020 => x"0c080000",
  2021 => x"0c060306",
  2022 => x"80800008",
  2023 => x"80808080",
  2024 => x"00000080",
  2025 => x"04070300",
  2026 => x"20000000",
  2027 => x"7c545474",
  2028 => x"7f000078",
  2029 => x"7c44447f",
  2030 => x"38000038",
  2031 => x"4444447c",
  2032 => x"38000000",
  2033 => x"7f44447c",
  2034 => x"3800007f",
  2035 => x"5c54547c",
  2036 => x"04000018",
  2037 => x"05057f7e",
  2038 => x"18000000",
  2039 => x"fca4a4bc",
  2040 => x"7f00007c",
  2041 => x"7c04047f",
  2042 => x"00000078",
  2043 => x"407d3d00",
  2044 => x"80000000",
  2045 => x"7dfd8080",
  2046 => x"7f000000",
  2047 => x"6c38107f",
  2048 => x"00000044",
  2049 => x"407f3f00",
  2050 => x"7c7c0000",
  2051 => x"7c0c180c",
  2052 => x"7c000078",
  2053 => x"7c04047c",
  2054 => x"38000078",
  2055 => x"7c44447c",
  2056 => x"fc000038",
  2057 => x"3c2424fc",
  2058 => x"18000018",
  2059 => x"fc24243c",
  2060 => x"7c0000fc",
  2061 => x"0c04047c",
  2062 => x"48000008",
  2063 => x"7454545c",
  2064 => x"04000020",
  2065 => x"44447f3f",
  2066 => x"3c000000",
  2067 => x"7c40407c",
  2068 => x"1c00007c",
  2069 => x"3c60603c",
  2070 => x"7c3c001c",
  2071 => x"7c603060",
  2072 => x"6c44003c",
  2073 => x"6c381038",
  2074 => x"1c000044",
  2075 => x"3c60e0bc",
  2076 => x"4400001c",
  2077 => x"4c5c7464",
  2078 => x"08000044",
  2079 => x"41773e08",
  2080 => x"00000041",
  2081 => x"007f7f00",
  2082 => x"41000000",
  2083 => x"083e7741",
  2084 => x"01020008",
  2085 => x"02020301",
  2086 => x"7f7f0001",
  2087 => x"7f7f7f7f",
  2088 => x"0808007f",
  2089 => x"3e3e1c1c",
  2090 => x"7f7f7f7f",
  2091 => x"1c1c3e3e",
  2092 => x"10000808",
  2093 => x"187c7c18",
  2094 => x"10000010",
  2095 => x"307c7c30",
  2096 => x"30100010",
  2097 => x"1e786060",
  2098 => x"66420006",
  2099 => x"663c183c",
  2100 => x"38780042",
  2101 => x"6cc6c26a",
  2102 => x"00600038",
  2103 => x"00006000",
  2104 => x"5e0e0060",
  2105 => x"0e5d5c5b",
  2106 => x"c24c711e",
  2107 => x"4dbffdec",
  2108 => x"1ec04bc0",
  2109 => x"c702ab74",
  2110 => x"48a6c487",
  2111 => x"87c578c0",
  2112 => x"c148a6c4",
  2113 => x"1e66c478",
  2114 => x"dfee4973",
  2115 => x"c086c887",
  2116 => x"eeef49e0",
  2117 => x"4aa5c487",
  2118 => x"f0f0496a",
  2119 => x"87c6f187",
  2120 => x"83c185cb",
  2121 => x"04abb7c8",
  2122 => x"2687c7ff",
  2123 => x"4c264d26",
  2124 => x"4f264b26",
  2125 => x"c24a711e",
  2126 => x"c25ac1ed",
  2127 => x"c748c1ed",
  2128 => x"ddfe4978",
  2129 => x"1e4f2687",
  2130 => x"4a711e73",
  2131 => x"03aab7c0",
  2132 => x"d3c287d3",
  2133 => x"c405bfc3",
  2134 => x"c24bc187",
  2135 => x"c24bc087",
  2136 => x"c45bc7d3",
  2137 => x"c7d3c287",
  2138 => x"c3d3c25a",
  2139 => x"9ac14abf",
  2140 => x"49a2c0c1",
  2141 => x"fc87e8ec",
  2142 => x"c3d3c248",
  2143 => x"effe78bf",
  2144 => x"4a711e87",
  2145 => x"721e66c4",
  2146 => x"87f9ea49",
  2147 => x"1e4f2626",
  2148 => x"c348d4ff",
  2149 => x"d0ff78ff",
  2150 => x"78e1c048",
  2151 => x"c148d4ff",
  2152 => x"c4487178",
  2153 => x"08d4ff30",
  2154 => x"48d0ff78",
  2155 => x"2678e0c0",
  2156 => x"d3c21e4f",
  2157 => x"e649bfc3",
  2158 => x"ecc287f9",
  2159 => x"bfe848f5",
  2160 => x"f1ecc278",
  2161 => x"78bfec48",
  2162 => x"bff5ecc2",
  2163 => x"ffc3494a",
  2164 => x"2ab7c899",
  2165 => x"b0714872",
  2166 => x"58fdecc2",
  2167 => x"5e0e4f26",
  2168 => x"0e5d5c5b",
  2169 => x"c8ff4b71",
  2170 => x"f0ecc287",
  2171 => x"7350c048",
  2172 => x"87dfe649",
  2173 => x"c24c4970",
  2174 => x"49eecb9c",
  2175 => x"7087cccb",
  2176 => x"f0ecc24d",
  2177 => x"c105bf97",
  2178 => x"66d087e2",
  2179 => x"f9ecc249",
  2180 => x"d60599bf",
  2181 => x"4966d487",
  2182 => x"bff1ecc2",
  2183 => x"87cb0599",
  2184 => x"eee54973",
  2185 => x"02987087",
  2186 => x"c187c1c1",
  2187 => x"87c1fe4c",
  2188 => x"e2ca4975",
  2189 => x"02987087",
  2190 => x"ecc287c6",
  2191 => x"50c148f0",
  2192 => x"97f0ecc2",
  2193 => x"e3c005bf",
  2194 => x"f9ecc287",
  2195 => x"66d049bf",
  2196 => x"d6ff0599",
  2197 => x"f1ecc287",
  2198 => x"66d449bf",
  2199 => x"caff0599",
  2200 => x"e4497387",
  2201 => x"987087ed",
  2202 => x"87fffe05",
  2203 => x"fbfa4874",
  2204 => x"5b5e0e87",
  2205 => x"f80e5d5c",
  2206 => x"4c4dc086",
  2207 => x"c47ebfec",
  2208 => x"ecc248a6",
  2209 => x"c178bffd",
  2210 => x"c71ec01e",
  2211 => x"87cefd49",
  2212 => x"987086c8",
  2213 => x"ff87cd02",
  2214 => x"87ebfa49",
  2215 => x"e349dac1",
  2216 => x"4dc187f1",
  2217 => x"97f0ecc2",
  2218 => x"87cf02bf",
  2219 => x"bffbd2c2",
  2220 => x"c2b9c149",
  2221 => x"7159ffd2",
  2222 => x"c287d4fb",
  2223 => x"4bbff5ec",
  2224 => x"bfc3d3c2",
  2225 => x"87e9c005",
  2226 => x"e349fdc3",
  2227 => x"fac387c5",
  2228 => x"87ffe249",
  2229 => x"ffc34973",
  2230 => x"c01e7199",
  2231 => x"87e1fa49",
  2232 => x"b7c84973",
  2233 => x"c11e7129",
  2234 => x"87d5fa49",
  2235 => x"f4c586c8",
  2236 => x"f9ecc287",
  2237 => x"029b4bbf",
  2238 => x"d2c287dd",
  2239 => x"c749bfff",
  2240 => x"987087d5",
  2241 => x"c087c405",
  2242 => x"c287d24b",
  2243 => x"fac649e0",
  2244 => x"c3d3c287",
  2245 => x"c287c658",
  2246 => x"c048ffd2",
  2247 => x"c2497378",
  2248 => x"87cd0599",
  2249 => x"e149ebc3",
  2250 => x"497087e9",
  2251 => x"c20299c2",
  2252 => x"734cfb87",
  2253 => x"0599c149",
  2254 => x"f4c387cd",
  2255 => x"87d3e149",
  2256 => x"99c24970",
  2257 => x"fa87c202",
  2258 => x"c849734c",
  2259 => x"87cd0599",
  2260 => x"e049f5c3",
  2261 => x"497087fd",
  2262 => x"d50299c2",
  2263 => x"c1edc287",
  2264 => x"87ca02bf",
  2265 => x"c288c148",
  2266 => x"c058c5ed",
  2267 => x"4cff87c2",
  2268 => x"49734dc1",
  2269 => x"cd0599c4",
  2270 => x"49f2c387",
  2271 => x"7087d4e0",
  2272 => x"0299c249",
  2273 => x"edc287dc",
  2274 => x"487ebfc1",
  2275 => x"03a8b7c7",
  2276 => x"6e87cbc0",
  2277 => x"c280c148",
  2278 => x"c058c5ed",
  2279 => x"4cfe87c2",
  2280 => x"fdc34dc1",
  2281 => x"eadfff49",
  2282 => x"c2497087",
  2283 => x"87d50299",
  2284 => x"bfc1edc2",
  2285 => x"87c9c002",
  2286 => x"48c1edc2",
  2287 => x"c2c078c0",
  2288 => x"c14cfd87",
  2289 => x"49fac34d",
  2290 => x"87c7dfff",
  2291 => x"99c24970",
  2292 => x"87d9c002",
  2293 => x"bfc1edc2",
  2294 => x"a8b7c748",
  2295 => x"87c9c003",
  2296 => x"48c1edc2",
  2297 => x"c2c078c7",
  2298 => x"c14cfc87",
  2299 => x"acb7c04d",
  2300 => x"87d3c003",
  2301 => x"c14866c4",
  2302 => x"7e7080d8",
  2303 => x"c002bf6e",
  2304 => x"744b87c5",
  2305 => x"c00f7349",
  2306 => x"1ef0c31e",
  2307 => x"f749dac1",
  2308 => x"86c887cc",
  2309 => x"c0029870",
  2310 => x"edc287d8",
  2311 => x"6e7ebfc1",
  2312 => x"c491cb49",
  2313 => x"82714a66",
  2314 => x"c5c0026a",
  2315 => x"496e4b87",
  2316 => x"9d750f73",
  2317 => x"87c8c002",
  2318 => x"bfc1edc2",
  2319 => x"87e2f249",
  2320 => x"bfc7d3c2",
  2321 => x"87ddc002",
  2322 => x"87cbc249",
  2323 => x"c0029870",
  2324 => x"edc287d3",
  2325 => x"f249bfc1",
  2326 => x"49c087c8",
  2327 => x"c287e8f3",
  2328 => x"c048c7d3",
  2329 => x"f38ef878",
  2330 => x"5e0e87c2",
  2331 => x"0e5d5c5b",
  2332 => x"c24c711e",
  2333 => x"49bffdec",
  2334 => x"4da1cdc1",
  2335 => x"6981d1c1",
  2336 => x"029c747e",
  2337 => x"a5c487cf",
  2338 => x"c27b744b",
  2339 => x"49bffdec",
  2340 => x"6e87e1f2",
  2341 => x"059c747b",
  2342 => x"4bc087c4",
  2343 => x"4bc187c2",
  2344 => x"e2f24973",
  2345 => x"0266d487",
  2346 => x"de4987c7",
  2347 => x"c24a7087",
  2348 => x"c24ac087",
  2349 => x"265acbd3",
  2350 => x"0087f1f1",
  2351 => x"00000000",
  2352 => x"00000000",
  2353 => x"00000000",
  2354 => x"1e000000",
  2355 => x"c8ff4a71",
  2356 => x"a17249bf",
  2357 => x"1e4f2648",
  2358 => x"89bfc8ff",
  2359 => x"c0c0c0fe",
  2360 => x"01a9c0c0",
  2361 => x"4ac087c4",
  2362 => x"4ac187c2",
  2363 => x"4f264872",
  2364 => x"5c5b5e0e",
  2365 => x"4b710e5d",
  2366 => x"d04cd4ff",
  2367 => x"78c04866",
  2368 => x"dcff49d6",
  2369 => x"ffc387c5",
  2370 => x"c3496c7c",
  2371 => x"4d7199ff",
  2372 => x"99f0c349",
  2373 => x"05a9e0c1",
  2374 => x"ffc387cb",
  2375 => x"c3486c7c",
  2376 => x"0866d098",
  2377 => x"7cffc378",
  2378 => x"c8494a6c",
  2379 => x"7cffc331",
  2380 => x"b2714a6c",
  2381 => x"31c84972",
  2382 => x"6c7cffc3",
  2383 => x"72b2714a",
  2384 => x"c331c849",
  2385 => x"4a6c7cff",
  2386 => x"d0ffb271",
  2387 => x"78e0c048",
  2388 => x"c2029b73",
  2389 => x"757b7287",
  2390 => x"264d2648",
  2391 => x"264b264c",
  2392 => x"4f261e4f",
  2393 => x"5c5b5e0e",
  2394 => x"7686f80e",
  2395 => x"49a6c81e",
  2396 => x"c487fdfd",
  2397 => x"6e4b7086",
  2398 => x"03a8c448",
  2399 => x"7387f0c2",
  2400 => x"9af0c34a",
  2401 => x"02aad0c1",
  2402 => x"e0c187c7",
  2403 => x"dec205aa",
  2404 => x"c8497387",
  2405 => x"87c30299",
  2406 => x"7387c6ff",
  2407 => x"c29cc34c",
  2408 => x"c2c105ac",
  2409 => x"4966c487",
  2410 => x"1e7131c9",
  2411 => x"d44a66c4",
  2412 => x"c5edc292",
  2413 => x"fe817249",
  2414 => x"d887ced0",
  2415 => x"cad9ff49",
  2416 => x"1ec0c887",
  2417 => x"49e2dbc2",
  2418 => x"87d2ecfd",
  2419 => x"c048d0ff",
  2420 => x"dbc278e0",
  2421 => x"66cc1ee2",
  2422 => x"c292d44a",
  2423 => x"7249c5ed",
  2424 => x"d6cefe81",
  2425 => x"c186cc87",
  2426 => x"c2c105ac",
  2427 => x"4966c487",
  2428 => x"1e7131c9",
  2429 => x"d44a66c4",
  2430 => x"c5edc292",
  2431 => x"fe817249",
  2432 => x"c287c6cf",
  2433 => x"c81ee2db",
  2434 => x"92d44a66",
  2435 => x"49c5edc2",
  2436 => x"ccfe8172",
  2437 => x"49d787d7",
  2438 => x"87efd7ff",
  2439 => x"c21ec0c8",
  2440 => x"fd49e2db",
  2441 => x"cc87d0ea",
  2442 => x"48d0ff86",
  2443 => x"f878e0c0",
  2444 => x"87e7fc8e",
  2445 => x"5c5b5e0e",
  2446 => x"711e0e5d",
  2447 => x"4cd4ff4d",
  2448 => x"487e66d4",
  2449 => x"06a8b7c3",
  2450 => x"48c087c5",
  2451 => x"7587e9c1",
  2452 => x"fedcfe49",
  2453 => x"c41e7587",
  2454 => x"93d44b66",
  2455 => x"83c5edc2",
  2456 => x"c6fe4973",
  2457 => x"83c887d3",
  2458 => x"d0ff4b6b",
  2459 => x"78e1c848",
  2460 => x"48737cdd",
  2461 => x"7098ffc3",
  2462 => x"c849737c",
  2463 => x"487129b7",
  2464 => x"7098ffc3",
  2465 => x"d049737c",
  2466 => x"487129b7",
  2467 => x"7098ffc3",
  2468 => x"d848737c",
  2469 => x"7c7028b7",
  2470 => x"7c7c7cc0",
  2471 => x"7c7c7c7c",
  2472 => x"7c7c7c7c",
  2473 => x"48d0ff7c",
  2474 => x"c478e0c0",
  2475 => x"49dc1e66",
  2476 => x"87fcd5ff",
  2477 => x"487386c8",
  2478 => x"87ddfa26",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
