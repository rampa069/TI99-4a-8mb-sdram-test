
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d8",x"ee",x"c2"),
    14 => (x"48",x"fc",x"da",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f4",x"e2"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"fc",x"da"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"da",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"fc"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"c0",x"db",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"c4",x"db",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"c4",x"db",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"c4",x"db"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"cb",x"db"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"cc",x"db"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"cd",x"db",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"db",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"cd"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"ce",x"db",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"c9",x"db"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"ca",x"db",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"db",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"cb"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"cc",x"db",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e3",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"ea"),
   330 => (x"1e",x"e2",x"db",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"e2",x"f2",x"c0",x"7e"),
   337 => (x"dc",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"d8"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"de",x"f2"),
   343 => (x"4a",x"f4",x"dc",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e2",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"e8"),
   350 => (x"bf",x"9f",x"e0",x"e3"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"e8",x"e2",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"db",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"e2"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"de",x"f2"),
   365 => (x"4a",x"f4",x"dc",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"ea",x"e3"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"e2",x"f2"),
   372 => (x"4a",x"d8",x"dc",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"e0",x"e3",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e3",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"e1"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"e2",x"db",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"ed",x"db",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"ee",x"db"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"ef",x"db",x"c2"),
   400 => (x"e3",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"e6"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"ea",x"e3"),
   404 => (x"bf",x"97",x"f0",x"db"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"f1",x"db"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e7",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"f7"),
   410 => (x"97",x"f2",x"db",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"ea",x"e3",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"de",x"f2",x"c0",x"87"),
   415 => (x"dc",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"f4"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"e2",x"e3"),
   422 => (x"5c",x"cb",x"e8",x"c2"),
   423 => (x"97",x"c7",x"dc",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"c6",x"dc",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"c8",x"dc",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"c9",x"dc"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"f7",x"e7",x"c2",x"91"),
   434 => (x"e7",x"c2",x"81",x"bf"),
   435 => (x"dc",x"c2",x"59",x"ff"),
   436 => (x"4a",x"bf",x"97",x"cf"),
   437 => (x"dc",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"ce"),
   439 => (x"dc",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"d0"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"d1",x"dc",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e8",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"c3"),
   447 => (x"e8",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"c3"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"f4",x"db",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"f3",x"db",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"cb",x"e8"),
   457 => (x"bf",x"97",x"f9",x"db"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"f8",x"db"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"c7",x"e8",x"c2"),
   463 => (x"48",x"ff",x"e7",x"c2"),
   464 => (x"e7",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"fb"),
   466 => (x"cb",x"e8",x"c2",x"78"),
   467 => (x"ff",x"e7",x"c2",x"48"),
   468 => (x"e8",x"c2",x"78",x"bf"),
   469 => (x"e8",x"c2",x"48",x"cf"),
   470 => (x"c2",x"78",x"bf",x"c3"),
   471 => (x"02",x"bf",x"ea",x"e3"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"c7",x"e8",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"ee",x"e3",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"ea",x"e3"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e7",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"f7"),
   492 => (x"ab",x"bf",x"da",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"de",x"f2"),
   495 => (x"73",x"1e",x"e2",x"db"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"ea",x"e3",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"e2",x"db"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"e2",x"db",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c1",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"ea",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d6",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"f2",x"e3",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d4",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"cf",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"ea",x"e3"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"49",x"6e",x"7e",x"c0"),
   556 => (x"bf",x"66",x"c4",x"48"),
   557 => (x"08",x"66",x"c4",x"80"),
   558 => (x"cc",x"7c",x"c0",x"78"),
   559 => (x"66",x"c4",x"49",x"a4"),
   560 => (x"a4",x"d0",x"79",x"bf"),
   561 => (x"c1",x"79",x"c0",x"49"),
   562 => (x"c0",x"87",x"c2",x"48"),
   563 => (x"fa",x"8e",x"f8",x"48"),
   564 => (x"5e",x"0e",x"87",x"ed"),
   565 => (x"0e",x"5d",x"5c",x"5b"),
   566 => (x"02",x"9c",x"4c",x"71"),
   567 => (x"c8",x"87",x"cb",x"c1"),
   568 => (x"02",x"69",x"49",x"a4"),
   569 => (x"d0",x"87",x"c3",x"c1"),
   570 => (x"49",x"6c",x"4a",x"66"),
   571 => (x"72",x"48",x"a6",x"d0"),
   572 => (x"b9",x"4d",x"78",x"a1"),
   573 => (x"bf",x"e6",x"e3",x"c2"),
   574 => (x"72",x"ba",x"ff",x"4a"),
   575 => (x"02",x"99",x"71",x"99"),
   576 => (x"c4",x"87",x"e4",x"c0"),
   577 => (x"49",x"6b",x"4b",x"a4"),
   578 => (x"70",x"87",x"fc",x"f9"),
   579 => (x"e2",x"e3",x"c2",x"7b"),
   580 => (x"81",x"6c",x"49",x"bf"),
   581 => (x"b9",x"75",x"7c",x"71"),
   582 => (x"bf",x"e6",x"e3",x"c2"),
   583 => (x"72",x"ba",x"ff",x"4a"),
   584 => (x"05",x"99",x"71",x"99"),
   585 => (x"d0",x"87",x"dc",x"ff"),
   586 => (x"d2",x"f9",x"7c",x"66"),
   587 => (x"1e",x"73",x"1e",x"87"),
   588 => (x"02",x"9b",x"4b",x"71"),
   589 => (x"a3",x"c8",x"87",x"c7"),
   590 => (x"c5",x"05",x"69",x"49"),
   591 => (x"c0",x"48",x"c0",x"87"),
   592 => (x"e7",x"c2",x"87",x"f6"),
   593 => (x"c4",x"49",x"bf",x"fb"),
   594 => (x"4a",x"6a",x"4a",x"a3"),
   595 => (x"e3",x"c2",x"8a",x"c2"),
   596 => (x"72",x"92",x"bf",x"e2"),
   597 => (x"e3",x"c2",x"49",x"a1"),
   598 => (x"6b",x"4a",x"bf",x"e6"),
   599 => (x"49",x"a1",x"72",x"9a"),
   600 => (x"59",x"de",x"f2",x"c0"),
   601 => (x"71",x"1e",x"66",x"c8"),
   602 => (x"c4",x"87",x"e4",x"ea"),
   603 => (x"05",x"98",x"70",x"86"),
   604 => (x"48",x"c0",x"87",x"c4"),
   605 => (x"48",x"c1",x"87",x"c2"),
   606 => (x"1e",x"87",x"c8",x"f8"),
   607 => (x"4b",x"71",x"1e",x"73"),
   608 => (x"87",x"c7",x"02",x"9b"),
   609 => (x"69",x"49",x"a3",x"c8"),
   610 => (x"c0",x"87",x"c5",x"05"),
   611 => (x"87",x"f6",x"c0",x"48"),
   612 => (x"bf",x"fb",x"e7",x"c2"),
   613 => (x"4a",x"a3",x"c4",x"49"),
   614 => (x"8a",x"c2",x"4a",x"6a"),
   615 => (x"bf",x"e2",x"e3",x"c2"),
   616 => (x"49",x"a1",x"72",x"92"),
   617 => (x"bf",x"e6",x"e3",x"c2"),
   618 => (x"72",x"9a",x"6b",x"4a"),
   619 => (x"f2",x"c0",x"49",x"a1"),
   620 => (x"66",x"c8",x"59",x"de"),
   621 => (x"cf",x"e6",x"71",x"1e"),
   622 => (x"70",x"86",x"c4",x"87"),
   623 => (x"87",x"c4",x"05",x"98"),
   624 => (x"87",x"c2",x"48",x"c0"),
   625 => (x"fa",x"f6",x"48",x"c1"),
   626 => (x"5b",x"5e",x"0e",x"87"),
   627 => (x"1e",x"0e",x"5d",x"5c"),
   628 => (x"66",x"d4",x"4b",x"71"),
   629 => (x"02",x"9b",x"73",x"4d"),
   630 => (x"c8",x"87",x"cc",x"c1"),
   631 => (x"02",x"69",x"49",x"a3"),
   632 => (x"d0",x"87",x"c4",x"c1"),
   633 => (x"e3",x"c2",x"4c",x"a3"),
   634 => (x"ff",x"49",x"bf",x"e6"),
   635 => (x"99",x"4a",x"6c",x"b9"),
   636 => (x"a9",x"66",x"d4",x"7e"),
   637 => (x"c0",x"87",x"cd",x"06"),
   638 => (x"a3",x"cc",x"7c",x"7b"),
   639 => (x"49",x"a3",x"c4",x"4a"),
   640 => (x"87",x"ca",x"79",x"6a"),
   641 => (x"c0",x"f8",x"49",x"72"),
   642 => (x"4d",x"66",x"d4",x"99"),
   643 => (x"49",x"75",x"8d",x"71"),
   644 => (x"1e",x"71",x"29",x"c9"),
   645 => (x"f9",x"fa",x"49",x"73"),
   646 => (x"e2",x"db",x"c2",x"87"),
   647 => (x"fc",x"49",x"73",x"1e"),
   648 => (x"86",x"c8",x"87",x"cb"),
   649 => (x"26",x"7c",x"66",x"d4"),
   650 => (x"1e",x"87",x"d4",x"f5"),
   651 => (x"4b",x"71",x"1e",x"73"),
   652 => (x"e4",x"c0",x"02",x"9b"),
   653 => (x"cf",x"e8",x"c2",x"87"),
   654 => (x"c2",x"4a",x"73",x"5b"),
   655 => (x"e2",x"e3",x"c2",x"8a"),
   656 => (x"c2",x"92",x"49",x"bf"),
   657 => (x"48",x"bf",x"fb",x"e7"),
   658 => (x"e8",x"c2",x"80",x"72"),
   659 => (x"48",x"71",x"58",x"d3"),
   660 => (x"e3",x"c2",x"30",x"c4"),
   661 => (x"ed",x"c0",x"58",x"f2"),
   662 => (x"cb",x"e8",x"c2",x"87"),
   663 => (x"ff",x"e7",x"c2",x"48"),
   664 => (x"e8",x"c2",x"78",x"bf"),
   665 => (x"e8",x"c2",x"48",x"cf"),
   666 => (x"c2",x"78",x"bf",x"c3"),
   667 => (x"02",x"bf",x"ea",x"e3"),
   668 => (x"e3",x"c2",x"87",x"c9"),
   669 => (x"c4",x"49",x"bf",x"e2"),
   670 => (x"c2",x"87",x"c7",x"31"),
   671 => (x"49",x"bf",x"c7",x"e8"),
   672 => (x"e3",x"c2",x"31",x"c4"),
   673 => (x"fa",x"f3",x"59",x"f2"),
   674 => (x"5b",x"5e",x"0e",x"87"),
   675 => (x"4a",x"71",x"0e",x"5c"),
   676 => (x"9a",x"72",x"4b",x"c0"),
   677 => (x"87",x"e1",x"c0",x"02"),
   678 => (x"9f",x"49",x"a2",x"da"),
   679 => (x"e3",x"c2",x"4b",x"69"),
   680 => (x"cf",x"02",x"bf",x"ea"),
   681 => (x"49",x"a2",x"d4",x"87"),
   682 => (x"4c",x"49",x"69",x"9f"),
   683 => (x"9c",x"ff",x"ff",x"c0"),
   684 => (x"87",x"c2",x"34",x"d0"),
   685 => (x"49",x"74",x"4c",x"c0"),
   686 => (x"fd",x"49",x"73",x"b3"),
   687 => (x"c0",x"f3",x"87",x"ed"),
   688 => (x"5b",x"5e",x"0e",x"87"),
   689 => (x"f4",x"0e",x"5d",x"5c"),
   690 => (x"c0",x"4a",x"71",x"86"),
   691 => (x"02",x"9a",x"72",x"7e"),
   692 => (x"db",x"c2",x"87",x"d8"),
   693 => (x"78",x"c0",x"48",x"de"),
   694 => (x"48",x"d6",x"db",x"c2"),
   695 => (x"bf",x"cf",x"e8",x"c2"),
   696 => (x"da",x"db",x"c2",x"78"),
   697 => (x"cb",x"e8",x"c2",x"48"),
   698 => (x"e3",x"c2",x"78",x"bf"),
   699 => (x"50",x"c0",x"48",x"ff"),
   700 => (x"bf",x"ee",x"e3",x"c2"),
   701 => (x"de",x"db",x"c2",x"49"),
   702 => (x"aa",x"71",x"4a",x"bf"),
   703 => (x"87",x"c9",x"c4",x"03"),
   704 => (x"99",x"cf",x"49",x"72"),
   705 => (x"87",x"e9",x"c0",x"05"),
   706 => (x"48",x"da",x"f2",x"c0"),
   707 => (x"bf",x"d6",x"db",x"c2"),
   708 => (x"e2",x"db",x"c2",x"78"),
   709 => (x"d6",x"db",x"c2",x"1e"),
   710 => (x"db",x"c2",x"49",x"bf"),
   711 => (x"a1",x"c1",x"48",x"d6"),
   712 => (x"ea",x"e3",x"71",x"78"),
   713 => (x"c0",x"86",x"c4",x"87"),
   714 => (x"c2",x"48",x"d6",x"f2"),
   715 => (x"cc",x"78",x"e2",x"db"),
   716 => (x"d6",x"f2",x"c0",x"87"),
   717 => (x"e0",x"c0",x"48",x"bf"),
   718 => (x"da",x"f2",x"c0",x"80"),
   719 => (x"de",x"db",x"c2",x"58"),
   720 => (x"80",x"c1",x"48",x"bf"),
   721 => (x"58",x"e2",x"db",x"c2"),
   722 => (x"00",x"0c",x"96",x"27"),
   723 => (x"bf",x"97",x"bf",x"00"),
   724 => (x"c2",x"02",x"9d",x"4d"),
   725 => (x"e5",x"c3",x"87",x"e3"),
   726 => (x"dc",x"c2",x"02",x"ad"),
   727 => (x"d6",x"f2",x"c0",x"87"),
   728 => (x"a3",x"cb",x"4b",x"bf"),
   729 => (x"cf",x"4c",x"11",x"49"),
   730 => (x"d2",x"c1",x"05",x"ac"),
   731 => (x"df",x"49",x"75",x"87"),
   732 => (x"cd",x"89",x"c1",x"99"),
   733 => (x"f2",x"e3",x"c2",x"91"),
   734 => (x"4a",x"a3",x"c1",x"81"),
   735 => (x"a3",x"c3",x"51",x"12"),
   736 => (x"c5",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"c7"),
   739 => (x"4a",x"a3",x"c9",x"51"),
   740 => (x"a3",x"ce",x"51",x"12"),
   741 => (x"d0",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"12",x"4a",x"a3",x"d2"),
   744 => (x"4a",x"a3",x"d4",x"51"),
   745 => (x"a3",x"d6",x"51",x"12"),
   746 => (x"d8",x"51",x"12",x"4a"),
   747 => (x"51",x"12",x"4a",x"a3"),
   748 => (x"12",x"4a",x"a3",x"dc"),
   749 => (x"4a",x"a3",x"de",x"51"),
   750 => (x"7e",x"c1",x"51",x"12"),
   751 => (x"74",x"87",x"fa",x"c0"),
   752 => (x"05",x"99",x"c8",x"49"),
   753 => (x"74",x"87",x"eb",x"c0"),
   754 => (x"05",x"99",x"d0",x"49"),
   755 => (x"66",x"dc",x"87",x"d1"),
   756 => (x"87",x"cb",x"c0",x"02"),
   757 => (x"66",x"dc",x"49",x"73"),
   758 => (x"02",x"98",x"70",x"0f"),
   759 => (x"6e",x"87",x"d3",x"c0"),
   760 => (x"87",x"c6",x"c0",x"05"),
   761 => (x"48",x"f2",x"e3",x"c2"),
   762 => (x"f2",x"c0",x"50",x"c0"),
   763 => (x"c2",x"48",x"bf",x"d6"),
   764 => (x"e3",x"c2",x"87",x"df"),
   765 => (x"50",x"c0",x"48",x"ff"),
   766 => (x"ee",x"e3",x"c2",x"7e"),
   767 => (x"db",x"c2",x"49",x"bf"),
   768 => (x"71",x"4a",x"bf",x"de"),
   769 => (x"f7",x"fb",x"04",x"aa"),
   770 => (x"cf",x"e8",x"c2",x"87"),
   771 => (x"c8",x"c0",x"05",x"bf"),
   772 => (x"ea",x"e3",x"c2",x"87"),
   773 => (x"f6",x"c1",x"02",x"bf"),
   774 => (x"da",x"db",x"c2",x"87"),
   775 => (x"e6",x"ed",x"49",x"bf"),
   776 => (x"de",x"db",x"c2",x"87"),
   777 => (x"48",x"a6",x"c4",x"58"),
   778 => (x"bf",x"da",x"db",x"c2"),
   779 => (x"ea",x"e3",x"c2",x"78"),
   780 => (x"d8",x"c0",x"02",x"bf"),
   781 => (x"49",x"66",x"c4",x"87"),
   782 => (x"ff",x"ff",x"ff",x"cf"),
   783 => (x"02",x"a9",x"99",x"f8"),
   784 => (x"c0",x"87",x"c5",x"c0"),
   785 => (x"87",x"e1",x"c0",x"4c"),
   786 => (x"dc",x"c0",x"4c",x"c1"),
   787 => (x"49",x"66",x"c4",x"87"),
   788 => (x"99",x"f8",x"ff",x"cf"),
   789 => (x"c8",x"c0",x"02",x"a9"),
   790 => (x"48",x"a6",x"c8",x"87"),
   791 => (x"c5",x"c0",x"78",x"c0"),
   792 => (x"48",x"a6",x"c8",x"87"),
   793 => (x"66",x"c8",x"78",x"c1"),
   794 => (x"05",x"9c",x"74",x"4c"),
   795 => (x"c4",x"87",x"e0",x"c0"),
   796 => (x"89",x"c2",x"49",x"66"),
   797 => (x"bf",x"e2",x"e3",x"c2"),
   798 => (x"e7",x"c2",x"91",x"4a"),
   799 => (x"c2",x"4a",x"bf",x"fb"),
   800 => (x"72",x"48",x"d6",x"db"),
   801 => (x"db",x"c2",x"78",x"a1"),
   802 => (x"78",x"c0",x"48",x"de"),
   803 => (x"c0",x"87",x"e1",x"f9"),
   804 => (x"eb",x"8e",x"f4",x"48"),
   805 => (x"00",x"00",x"87",x"e9"),
   806 => (x"ff",x"ff",x"00",x"00"),
   807 => (x"0c",x"a6",x"ff",x"ff"),
   808 => (x"0c",x"af",x"00",x"00"),
   809 => (x"41",x"46",x"00",x"00"),
   810 => (x"20",x"32",x"33",x"54"),
   811 => (x"46",x"00",x"20",x"20"),
   812 => (x"36",x"31",x"54",x"41"),
   813 => (x"00",x"20",x"20",x"20"),
   814 => (x"48",x"d4",x"ff",x"1e"),
   815 => (x"68",x"78",x"ff",x"c3"),
   816 => (x"1e",x"4f",x"26",x"48"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"d0",x"ff",x"78",x"ff"),
   819 => (x"78",x"e1",x"c0",x"48"),
   820 => (x"d4",x"48",x"d4",x"ff"),
   821 => (x"d3",x"e8",x"c2",x"78"),
   822 => (x"bf",x"d4",x"ff",x"48"),
   823 => (x"1e",x"4f",x"26",x"50"),
   824 => (x"c0",x"48",x"d0",x"ff"),
   825 => (x"4f",x"26",x"78",x"e0"),
   826 => (x"87",x"cc",x"ff",x"1e"),
   827 => (x"02",x"99",x"49",x"70"),
   828 => (x"fb",x"c0",x"87",x"c6"),
   829 => (x"87",x"f1",x"05",x"a9"),
   830 => (x"4f",x"26",x"48",x"71"),
   831 => (x"5c",x"5b",x"5e",x"0e"),
   832 => (x"c0",x"4b",x"71",x"0e"),
   833 => (x"87",x"f0",x"fe",x"4c"),
   834 => (x"02",x"99",x"49",x"70"),
   835 => (x"c0",x"87",x"f9",x"c0"),
   836 => (x"c0",x"02",x"a9",x"ec"),
   837 => (x"fb",x"c0",x"87",x"f2"),
   838 => (x"eb",x"c0",x"02",x"a9"),
   839 => (x"b7",x"66",x"cc",x"87"),
   840 => (x"87",x"c7",x"03",x"ac"),
   841 => (x"c2",x"02",x"66",x"d0"),
   842 => (x"71",x"53",x"71",x"87"),
   843 => (x"87",x"c2",x"02",x"99"),
   844 => (x"c3",x"fe",x"84",x"c1"),
   845 => (x"99",x"49",x"70",x"87"),
   846 => (x"c0",x"87",x"cd",x"02"),
   847 => (x"c7",x"02",x"a9",x"ec"),
   848 => (x"a9",x"fb",x"c0",x"87"),
   849 => (x"87",x"d5",x"ff",x"05"),
   850 => (x"c3",x"02",x"66",x"d0"),
   851 => (x"7b",x"97",x"c0",x"87"),
   852 => (x"05",x"a9",x"ec",x"c0"),
   853 => (x"4a",x"74",x"87",x"c4"),
   854 => (x"4a",x"74",x"87",x"c5"),
   855 => (x"72",x"8a",x"0a",x"c0"),
   856 => (x"26",x"87",x"c2",x"48"),
   857 => (x"26",x"4c",x"26",x"4d"),
   858 => (x"1e",x"4f",x"26",x"4b"),
   859 => (x"70",x"87",x"c9",x"fd"),
   860 => (x"aa",x"f0",x"c0",x"4a"),
   861 => (x"c0",x"87",x"c9",x"04"),
   862 => (x"c3",x"01",x"aa",x"f9"),
   863 => (x"8a",x"f0",x"c0",x"87"),
   864 => (x"04",x"aa",x"c1",x"c1"),
   865 => (x"da",x"c1",x"87",x"c9"),
   866 => (x"87",x"c3",x"01",x"aa"),
   867 => (x"72",x"8a",x"f7",x"c0"),
   868 => (x"0e",x"4f",x"26",x"48"),
   869 => (x"0e",x"5c",x"5b",x"5e"),
   870 => (x"d4",x"ff",x"4a",x"71"),
   871 => (x"c0",x"49",x"72",x"4b"),
   872 => (x"4c",x"70",x"87",x"e7"),
   873 => (x"87",x"c2",x"02",x"9c"),
   874 => (x"d0",x"ff",x"8c",x"c1"),
   875 => (x"c1",x"78",x"c5",x"48"),
   876 => (x"49",x"74",x"7b",x"d5"),
   877 => (x"e4",x"c1",x"31",x"c6"),
   878 => (x"4a",x"bf",x"97",x"d5"),
   879 => (x"70",x"b0",x"71",x"48"),
   880 => (x"48",x"d0",x"ff",x"7b"),
   881 => (x"dc",x"fe",x"78",x"c4"),
   882 => (x"5b",x"5e",x"0e",x"87"),
   883 => (x"f8",x"0e",x"5d",x"5c"),
   884 => (x"c0",x"4c",x"71",x"86"),
   885 => (x"87",x"eb",x"fb",x"7e"),
   886 => (x"f9",x"c0",x"4b",x"c0"),
   887 => (x"49",x"bf",x"97",x"f6"),
   888 => (x"cf",x"04",x"a9",x"c0"),
   889 => (x"87",x"c0",x"fc",x"87"),
   890 => (x"f9",x"c0",x"83",x"c1"),
   891 => (x"49",x"bf",x"97",x"f6"),
   892 => (x"87",x"f1",x"06",x"ab"),
   893 => (x"97",x"f6",x"f9",x"c0"),
   894 => (x"87",x"cf",x"02",x"bf"),
   895 => (x"70",x"87",x"f9",x"fa"),
   896 => (x"c6",x"02",x"99",x"49"),
   897 => (x"a9",x"ec",x"c0",x"87"),
   898 => (x"c0",x"87",x"f1",x"05"),
   899 => (x"87",x"e8",x"fa",x"4b"),
   900 => (x"e3",x"fa",x"4d",x"70"),
   901 => (x"58",x"a6",x"c8",x"87"),
   902 => (x"70",x"87",x"dd",x"fa"),
   903 => (x"c8",x"83",x"c1",x"4a"),
   904 => (x"69",x"97",x"49",x"a4"),
   905 => (x"c7",x"02",x"ad",x"49"),
   906 => (x"ad",x"ff",x"c0",x"87"),
   907 => (x"87",x"e7",x"c0",x"05"),
   908 => (x"97",x"49",x"a4",x"c9"),
   909 => (x"66",x"c4",x"49",x"69"),
   910 => (x"87",x"c7",x"02",x"a9"),
   911 => (x"a8",x"ff",x"c0",x"48"),
   912 => (x"ca",x"87",x"d4",x"05"),
   913 => (x"69",x"97",x"49",x"a4"),
   914 => (x"c6",x"02",x"aa",x"49"),
   915 => (x"aa",x"ff",x"c0",x"87"),
   916 => (x"c1",x"87",x"c4",x"05"),
   917 => (x"c0",x"87",x"d0",x"7e"),
   918 => (x"c6",x"02",x"ad",x"ec"),
   919 => (x"ad",x"fb",x"c0",x"87"),
   920 => (x"c0",x"87",x"c4",x"05"),
   921 => (x"6e",x"7e",x"c1",x"4b"),
   922 => (x"87",x"e1",x"fe",x"02"),
   923 => (x"73",x"87",x"f0",x"f9"),
   924 => (x"fb",x"8e",x"f8",x"48"),
   925 => (x"0e",x"00",x"87",x"ed"),
   926 => (x"5d",x"5c",x"5b",x"5e"),
   927 => (x"71",x"86",x"f8",x"0e"),
   928 => (x"4b",x"d4",x"ff",x"4d"),
   929 => (x"e8",x"c2",x"1e",x"75"),
   930 => (x"ec",x"e5",x"49",x"d8"),
   931 => (x"70",x"86",x"c4",x"87"),
   932 => (x"ca",x"c4",x"02",x"98"),
   933 => (x"48",x"a6",x"c4",x"87"),
   934 => (x"bf",x"d7",x"e4",x"c1"),
   935 => (x"fb",x"49",x"75",x"78"),
   936 => (x"d0",x"ff",x"87",x"f1"),
   937 => (x"c1",x"78",x"c5",x"48"),
   938 => (x"4a",x"c0",x"7b",x"d6"),
   939 => (x"11",x"49",x"a2",x"75"),
   940 => (x"cb",x"82",x"c1",x"7b"),
   941 => (x"f3",x"04",x"aa",x"b7"),
   942 => (x"c3",x"4a",x"cc",x"87"),
   943 => (x"82",x"c1",x"7b",x"ff"),
   944 => (x"aa",x"b7",x"e0",x"c0"),
   945 => (x"ff",x"87",x"f4",x"04"),
   946 => (x"78",x"c4",x"48",x"d0"),
   947 => (x"c5",x"7b",x"ff",x"c3"),
   948 => (x"7b",x"d3",x"c1",x"78"),
   949 => (x"78",x"c4",x"7b",x"c1"),
   950 => (x"b7",x"c0",x"48",x"66"),
   951 => (x"ee",x"c2",x"06",x"a8"),
   952 => (x"e0",x"e8",x"c2",x"87"),
   953 => (x"66",x"c4",x"4c",x"bf"),
   954 => (x"c8",x"88",x"74",x"48"),
   955 => (x"9c",x"74",x"58",x"a6"),
   956 => (x"87",x"f7",x"c1",x"02"),
   957 => (x"7e",x"e2",x"db",x"c2"),
   958 => (x"8c",x"4d",x"c0",x"c8"),
   959 => (x"03",x"ac",x"b7",x"c0"),
   960 => (x"c0",x"c8",x"87",x"c6"),
   961 => (x"4c",x"c0",x"4d",x"a4"),
   962 => (x"97",x"d3",x"e8",x"c2"),
   963 => (x"99",x"d0",x"49",x"bf"),
   964 => (x"c0",x"87",x"d0",x"02"),
   965 => (x"d8",x"e8",x"c2",x"1e"),
   966 => (x"87",x"d1",x"e8",x"49"),
   967 => (x"4a",x"70",x"86",x"c4"),
   968 => (x"c2",x"87",x"ed",x"c0"),
   969 => (x"c2",x"1e",x"e2",x"db"),
   970 => (x"e7",x"49",x"d8",x"e8"),
   971 => (x"86",x"c4",x"87",x"ff"),
   972 => (x"d0",x"ff",x"4a",x"70"),
   973 => (x"78",x"c5",x"c8",x"48"),
   974 => (x"6e",x"7b",x"d4",x"c1"),
   975 => (x"6e",x"7b",x"bf",x"97"),
   976 => (x"70",x"80",x"c1",x"48"),
   977 => (x"05",x"8d",x"c1",x"7e"),
   978 => (x"ff",x"87",x"f0",x"ff"),
   979 => (x"78",x"c4",x"48",x"d0"),
   980 => (x"c5",x"05",x"9a",x"72"),
   981 => (x"c1",x"48",x"c0",x"87"),
   982 => (x"1e",x"c1",x"87",x"c7"),
   983 => (x"49",x"d8",x"e8",x"c2"),
   984 => (x"c4",x"87",x"ef",x"e5"),
   985 => (x"05",x"9c",x"74",x"86"),
   986 => (x"c4",x"87",x"c9",x"fe"),
   987 => (x"b7",x"c0",x"48",x"66"),
   988 => (x"87",x"d1",x"06",x"a8"),
   989 => (x"48",x"d8",x"e8",x"c2"),
   990 => (x"80",x"d0",x"78",x"c0"),
   991 => (x"80",x"f4",x"78",x"c0"),
   992 => (x"bf",x"e4",x"e8",x"c2"),
   993 => (x"48",x"66",x"c4",x"78"),
   994 => (x"01",x"a8",x"b7",x"c0"),
   995 => (x"ff",x"87",x"d2",x"fd"),
   996 => (x"78",x"c5",x"48",x"d0"),
   997 => (x"c0",x"7b",x"d3",x"c1"),
   998 => (x"c1",x"78",x"c4",x"7b"),
   999 => (x"c0",x"87",x"c2",x"48"),
  1000 => (x"26",x"8e",x"f8",x"48"),
  1001 => (x"26",x"4c",x"26",x"4d"),
  1002 => (x"0e",x"4f",x"26",x"4b"),
  1003 => (x"5d",x"5c",x"5b",x"5e"),
  1004 => (x"4b",x"71",x"1e",x"0e"),
  1005 => (x"ab",x"4d",x"4c",x"c0"),
  1006 => (x"87",x"e8",x"c0",x"04"),
  1007 => (x"1e",x"c9",x"f7",x"c0"),
  1008 => (x"c4",x"02",x"9d",x"75"),
  1009 => (x"c2",x"4a",x"c0",x"87"),
  1010 => (x"72",x"4a",x"c1",x"87"),
  1011 => (x"87",x"f1",x"eb",x"49"),
  1012 => (x"7e",x"70",x"86",x"c4"),
  1013 => (x"05",x"6e",x"84",x"c1"),
  1014 => (x"4c",x"73",x"87",x"c2"),
  1015 => (x"ac",x"73",x"85",x"c1"),
  1016 => (x"87",x"d8",x"ff",x"06"),
  1017 => (x"fe",x"26",x"48",x"6e"),
  1018 => (x"5e",x"0e",x"87",x"f9"),
  1019 => (x"71",x"0e",x"5c",x"5b"),
  1020 => (x"02",x"66",x"cc",x"4b"),
  1021 => (x"c0",x"4c",x"87",x"d8"),
  1022 => (x"d8",x"02",x"8c",x"f0"),
  1023 => (x"c1",x"4a",x"74",x"87"),
  1024 => (x"87",x"d1",x"02",x"8a"),
  1025 => (x"87",x"cd",x"02",x"8a"),
  1026 => (x"87",x"c9",x"02",x"8a"),
  1027 => (x"49",x"73",x"87",x"d9"),
  1028 => (x"d2",x"87",x"e4",x"f9"),
  1029 => (x"c0",x"1e",x"74",x"87"),
  1030 => (x"d7",x"d8",x"c1",x"49"),
  1031 => (x"73",x"1e",x"74",x"87"),
  1032 => (x"cf",x"d8",x"c1",x"49"),
  1033 => (x"fd",x"86",x"c8",x"87"),
  1034 => (x"5e",x"0e",x"87",x"fb"),
  1035 => (x"0e",x"5d",x"5c",x"5b"),
  1036 => (x"49",x"4c",x"71",x"1e"),
  1037 => (x"e9",x"c2",x"91",x"de"),
  1038 => (x"85",x"71",x"4d",x"c0"),
  1039 => (x"c1",x"02",x"6d",x"97"),
  1040 => (x"e8",x"c2",x"87",x"dc"),
  1041 => (x"74",x"49",x"bf",x"ec"),
  1042 => (x"de",x"fd",x"71",x"81"),
  1043 => (x"48",x"7e",x"70",x"87"),
  1044 => (x"f2",x"c0",x"02",x"98"),
  1045 => (x"f4",x"e8",x"c2",x"87"),
  1046 => (x"cb",x"4a",x"70",x"4b"),
  1047 => (x"c6",x"c1",x"ff",x"49"),
  1048 => (x"cb",x"4b",x"74",x"87"),
  1049 => (x"e9",x"e4",x"c1",x"93"),
  1050 => (x"c1",x"83",x"c4",x"83"),
  1051 => (x"74",x"7b",x"e2",x"c2"),
  1052 => (x"ed",x"c1",x"c1",x"49"),
  1053 => (x"c1",x"7b",x"75",x"87"),
  1054 => (x"bf",x"97",x"d6",x"e4"),
  1055 => (x"e8",x"c2",x"1e",x"49"),
  1056 => (x"e5",x"fd",x"49",x"f4"),
  1057 => (x"74",x"86",x"c4",x"87"),
  1058 => (x"d5",x"c1",x"c1",x"49"),
  1059 => (x"c1",x"49",x"c0",x"87"),
  1060 => (x"c2",x"87",x"f4",x"c2"),
  1061 => (x"c0",x"48",x"d4",x"e8"),
  1062 => (x"dd",x"49",x"c1",x"78"),
  1063 => (x"fc",x"26",x"87",x"fb"),
  1064 => (x"6f",x"4c",x"87",x"c1"),
  1065 => (x"6e",x"69",x"64",x"61"),
  1066 => (x"2e",x"2e",x"2e",x"67"),
  1067 => (x"1e",x"73",x"1e",x"00"),
  1068 => (x"c2",x"49",x"4a",x"71"),
  1069 => (x"81",x"bf",x"ec",x"e8"),
  1070 => (x"87",x"ef",x"fb",x"71"),
  1071 => (x"02",x"9b",x"4b",x"70"),
  1072 => (x"e7",x"49",x"87",x"c4"),
  1073 => (x"e8",x"c2",x"87",x"c3"),
  1074 => (x"78",x"c0",x"48",x"ec"),
  1075 => (x"c8",x"dd",x"49",x"c1"),
  1076 => (x"87",x"d3",x"fb",x"87"),
  1077 => (x"c1",x"49",x"c0",x"1e"),
  1078 => (x"26",x"87",x"ec",x"c1"),
  1079 => (x"4a",x"71",x"1e",x"4f"),
  1080 => (x"c1",x"91",x"cb",x"49"),
  1081 => (x"c8",x"81",x"e9",x"e4"),
  1082 => (x"c2",x"48",x"11",x"81"),
  1083 => (x"c2",x"58",x"d8",x"e8"),
  1084 => (x"c0",x"48",x"ec",x"e8"),
  1085 => (x"dc",x"49",x"c1",x"78"),
  1086 => (x"4f",x"26",x"87",x"df"),
  1087 => (x"02",x"99",x"71",x"1e"),
  1088 => (x"e5",x"c1",x"87",x"d2"),
  1089 => (x"50",x"c0",x"48",x"fe"),
  1090 => (x"c3",x"c1",x"80",x"f7"),
  1091 => (x"e4",x"c1",x"40",x"dd"),
  1092 => (x"87",x"ce",x"78",x"e2"),
  1093 => (x"48",x"fa",x"e5",x"c1"),
  1094 => (x"78",x"db",x"e4",x"c1"),
  1095 => (x"c3",x"c1",x"80",x"fc"),
  1096 => (x"4f",x"26",x"78",x"d4"),
  1097 => (x"5c",x"5b",x"5e",x"0e"),
  1098 => (x"86",x"f4",x"0e",x"5d"),
  1099 => (x"4d",x"e2",x"db",x"c2"),
  1100 => (x"a6",x"c4",x"4c",x"c0"),
  1101 => (x"c2",x"78",x"c0",x"48"),
  1102 => (x"48",x"bf",x"ec",x"e8"),
  1103 => (x"c1",x"06",x"a8",x"c0"),
  1104 => (x"db",x"c2",x"87",x"c0"),
  1105 => (x"02",x"98",x"48",x"e2"),
  1106 => (x"c0",x"87",x"f7",x"c0"),
  1107 => (x"c8",x"1e",x"c9",x"f7"),
  1108 => (x"87",x"c7",x"02",x"66"),
  1109 => (x"c0",x"48",x"a6",x"c4"),
  1110 => (x"c4",x"87",x"c5",x"78"),
  1111 => (x"78",x"c1",x"48",x"a6"),
  1112 => (x"e5",x"49",x"66",x"c4"),
  1113 => (x"86",x"c4",x"87",x"db"),
  1114 => (x"84",x"c1",x"4d",x"70"),
  1115 => (x"c1",x"48",x"66",x"c4"),
  1116 => (x"58",x"a6",x"c8",x"80"),
  1117 => (x"bf",x"ec",x"e8",x"c2"),
  1118 => (x"87",x"c6",x"03",x"ac"),
  1119 => (x"ff",x"05",x"9d",x"75"),
  1120 => (x"4c",x"c0",x"87",x"c9"),
  1121 => (x"c3",x"02",x"9d",x"75"),
  1122 => (x"f7",x"c0",x"87",x"dc"),
  1123 => (x"66",x"c8",x"1e",x"c9"),
  1124 => (x"cc",x"87",x"c7",x"02"),
  1125 => (x"78",x"c0",x"48",x"a6"),
  1126 => (x"a6",x"cc",x"87",x"c5"),
  1127 => (x"cc",x"78",x"c1",x"48"),
  1128 => (x"dc",x"e4",x"49",x"66"),
  1129 => (x"70",x"86",x"c4",x"87"),
  1130 => (x"02",x"98",x"48",x"7e"),
  1131 => (x"49",x"87",x"e4",x"c2"),
  1132 => (x"69",x"97",x"81",x"cb"),
  1133 => (x"02",x"99",x"d0",x"49"),
  1134 => (x"74",x"87",x"d4",x"c1"),
  1135 => (x"c1",x"91",x"cb",x"49"),
  1136 => (x"c1",x"81",x"e9",x"e4"),
  1137 => (x"c8",x"79",x"ed",x"c2"),
  1138 => (x"51",x"ff",x"c3",x"81"),
  1139 => (x"91",x"de",x"49",x"74"),
  1140 => (x"4d",x"c0",x"e9",x"c2"),
  1141 => (x"c1",x"c2",x"85",x"71"),
  1142 => (x"a5",x"c1",x"7d",x"97"),
  1143 => (x"51",x"e0",x"c0",x"49"),
  1144 => (x"97",x"f2",x"e3",x"c2"),
  1145 => (x"87",x"d2",x"02",x"bf"),
  1146 => (x"a5",x"c2",x"84",x"c1"),
  1147 => (x"f2",x"e3",x"c2",x"4b"),
  1148 => (x"fe",x"49",x"db",x"4a"),
  1149 => (x"c1",x"87",x"f0",x"fa"),
  1150 => (x"a5",x"cd",x"87",x"d9"),
  1151 => (x"c1",x"51",x"c0",x"49"),
  1152 => (x"4b",x"a5",x"c2",x"84"),
  1153 => (x"49",x"cb",x"4a",x"6e"),
  1154 => (x"87",x"db",x"fa",x"fe"),
  1155 => (x"74",x"87",x"c4",x"c1"),
  1156 => (x"c1",x"91",x"cb",x"49"),
  1157 => (x"c1",x"81",x"e9",x"e4"),
  1158 => (x"c2",x"79",x"ea",x"c0"),
  1159 => (x"bf",x"97",x"f2",x"e3"),
  1160 => (x"74",x"87",x"d8",x"02"),
  1161 => (x"c1",x"91",x"de",x"49"),
  1162 => (x"c0",x"e9",x"c2",x"84"),
  1163 => (x"c2",x"83",x"71",x"4b"),
  1164 => (x"dd",x"4a",x"f2",x"e3"),
  1165 => (x"ee",x"f9",x"fe",x"49"),
  1166 => (x"74",x"87",x"d8",x"87"),
  1167 => (x"c2",x"93",x"de",x"4b"),
  1168 => (x"cb",x"83",x"c0",x"e9"),
  1169 => (x"51",x"c0",x"49",x"a3"),
  1170 => (x"6e",x"73",x"84",x"c1"),
  1171 => (x"fe",x"49",x"cb",x"4a"),
  1172 => (x"c4",x"87",x"d4",x"f9"),
  1173 => (x"80",x"c1",x"48",x"66"),
  1174 => (x"c7",x"58",x"a6",x"c8"),
  1175 => (x"c5",x"c0",x"03",x"ac"),
  1176 => (x"fc",x"05",x"6e",x"87"),
  1177 => (x"48",x"74",x"87",x"e4"),
  1178 => (x"f6",x"f4",x"8e",x"f4"),
  1179 => (x"1e",x"73",x"1e",x"87"),
  1180 => (x"cb",x"49",x"4b",x"71"),
  1181 => (x"e9",x"e4",x"c1",x"91"),
  1182 => (x"4a",x"a1",x"c8",x"81"),
  1183 => (x"48",x"d5",x"e4",x"c1"),
  1184 => (x"a1",x"c9",x"50",x"12"),
  1185 => (x"f6",x"f9",x"c0",x"4a"),
  1186 => (x"ca",x"50",x"12",x"48"),
  1187 => (x"d6",x"e4",x"c1",x"81"),
  1188 => (x"c1",x"50",x"11",x"48"),
  1189 => (x"bf",x"97",x"d6",x"e4"),
  1190 => (x"49",x"c0",x"1e",x"49"),
  1191 => (x"c2",x"87",x"cb",x"f5"),
  1192 => (x"de",x"48",x"d4",x"e8"),
  1193 => (x"d5",x"49",x"c1",x"78"),
  1194 => (x"f3",x"26",x"87",x"ef"),
  1195 => (x"5e",x"0e",x"87",x"f9"),
  1196 => (x"0e",x"5d",x"5c",x"5b"),
  1197 => (x"4d",x"71",x"86",x"f4"),
  1198 => (x"c1",x"91",x"cb",x"49"),
  1199 => (x"c8",x"81",x"e9",x"e4"),
  1200 => (x"a1",x"ca",x"4a",x"a1"),
  1201 => (x"48",x"a6",x"c4",x"7e"),
  1202 => (x"bf",x"dc",x"ec",x"c2"),
  1203 => (x"bf",x"97",x"6e",x"78"),
  1204 => (x"4c",x"66",x"c4",x"4b"),
  1205 => (x"48",x"12",x"2c",x"73"),
  1206 => (x"70",x"58",x"a6",x"cc"),
  1207 => (x"c9",x"84",x"c1",x"9c"),
  1208 => (x"49",x"69",x"97",x"81"),
  1209 => (x"c2",x"04",x"ac",x"b7"),
  1210 => (x"6e",x"4c",x"c0",x"87"),
  1211 => (x"c8",x"4a",x"bf",x"97"),
  1212 => (x"31",x"72",x"49",x"66"),
  1213 => (x"66",x"c4",x"b9",x"ff"),
  1214 => (x"72",x"48",x"74",x"99"),
  1215 => (x"48",x"4a",x"70",x"30"),
  1216 => (x"ec",x"c2",x"b0",x"71"),
  1217 => (x"e5",x"c0",x"58",x"e0"),
  1218 => (x"49",x"c0",x"87",x"d8"),
  1219 => (x"75",x"87",x"ca",x"d4"),
  1220 => (x"cd",x"f7",x"c0",x"49"),
  1221 => (x"f2",x"8e",x"f4",x"87"),
  1222 => (x"73",x"1e",x"87",x"c9"),
  1223 => (x"49",x"4b",x"71",x"1e"),
  1224 => (x"73",x"87",x"cb",x"fe"),
  1225 => (x"87",x"c6",x"fe",x"49"),
  1226 => (x"1e",x"87",x"fc",x"f1"),
  1227 => (x"4b",x"71",x"1e",x"73"),
  1228 => (x"02",x"4a",x"a3",x"c6"),
  1229 => (x"8a",x"c1",x"87",x"db"),
  1230 => (x"8a",x"87",x"d6",x"02"),
  1231 => (x"87",x"da",x"c1",x"02"),
  1232 => (x"fc",x"c0",x"02",x"8a"),
  1233 => (x"c0",x"02",x"8a",x"87"),
  1234 => (x"02",x"8a",x"87",x"e1"),
  1235 => (x"db",x"c1",x"87",x"cb"),
  1236 => (x"f6",x"49",x"c7",x"87"),
  1237 => (x"de",x"c1",x"87",x"c7"),
  1238 => (x"ec",x"e8",x"c2",x"87"),
  1239 => (x"cb",x"c1",x"02",x"bf"),
  1240 => (x"88",x"c1",x"48",x"87"),
  1241 => (x"58",x"f0",x"e8",x"c2"),
  1242 => (x"c2",x"87",x"c1",x"c1"),
  1243 => (x"02",x"bf",x"f0",x"e8"),
  1244 => (x"c2",x"87",x"f9",x"c0"),
  1245 => (x"48",x"bf",x"ec",x"e8"),
  1246 => (x"e8",x"c2",x"80",x"c1"),
  1247 => (x"eb",x"c0",x"58",x"f0"),
  1248 => (x"ec",x"e8",x"c2",x"87"),
  1249 => (x"89",x"c6",x"49",x"bf"),
  1250 => (x"59",x"f0",x"e8",x"c2"),
  1251 => (x"03",x"a9",x"b7",x"c0"),
  1252 => (x"e8",x"c2",x"87",x"da"),
  1253 => (x"78",x"c0",x"48",x"ec"),
  1254 => (x"e8",x"c2",x"87",x"d2"),
  1255 => (x"cb",x"02",x"bf",x"f0"),
  1256 => (x"ec",x"e8",x"c2",x"87"),
  1257 => (x"80",x"c6",x"48",x"bf"),
  1258 => (x"58",x"f0",x"e8",x"c2"),
  1259 => (x"e8",x"d1",x"49",x"c0"),
  1260 => (x"c0",x"49",x"73",x"87"),
  1261 => (x"ef",x"87",x"eb",x"f4"),
  1262 => (x"5e",x"0e",x"87",x"ed"),
  1263 => (x"0e",x"5d",x"5c",x"5b"),
  1264 => (x"dc",x"86",x"d4",x"ff"),
  1265 => (x"a6",x"c8",x"59",x"a6"),
  1266 => (x"c4",x"78",x"c0",x"48"),
  1267 => (x"66",x"c0",x"c1",x"80"),
  1268 => (x"c1",x"80",x"c4",x"78"),
  1269 => (x"c1",x"80",x"c4",x"78"),
  1270 => (x"f0",x"e8",x"c2",x"78"),
  1271 => (x"c2",x"78",x"c1",x"48"),
  1272 => (x"48",x"bf",x"d4",x"e8"),
  1273 => (x"c9",x"05",x"a8",x"de"),
  1274 => (x"87",x"f8",x"f4",x"87"),
  1275 => (x"cf",x"58",x"a6",x"cc"),
  1276 => (x"ce",x"e3",x"87",x"e6"),
  1277 => (x"87",x"f0",x"e3",x"87"),
  1278 => (x"70",x"87",x"fd",x"e2"),
  1279 => (x"ac",x"fb",x"c0",x"4c"),
  1280 => (x"87",x"fb",x"c1",x"02"),
  1281 => (x"c1",x"05",x"66",x"d8"),
  1282 => (x"fc",x"c0",x"87",x"ed"),
  1283 => (x"82",x"c4",x"4a",x"66"),
  1284 => (x"1e",x"72",x"7e",x"6a"),
  1285 => (x"48",x"cd",x"e0",x"c1"),
  1286 => (x"c8",x"49",x"66",x"c4"),
  1287 => (x"41",x"20",x"4a",x"a1"),
  1288 => (x"f9",x"05",x"aa",x"71"),
  1289 => (x"26",x"51",x"10",x"87"),
  1290 => (x"66",x"fc",x"c0",x"4a"),
  1291 => (x"ed",x"c9",x"c1",x"48"),
  1292 => (x"c7",x"49",x"6a",x"78"),
  1293 => (x"c0",x"51",x"74",x"81"),
  1294 => (x"c8",x"49",x"66",x"fc"),
  1295 => (x"c0",x"51",x"c1",x"81"),
  1296 => (x"c9",x"49",x"66",x"fc"),
  1297 => (x"c0",x"51",x"c0",x"81"),
  1298 => (x"ca",x"49",x"66",x"fc"),
  1299 => (x"c1",x"51",x"c0",x"81"),
  1300 => (x"6a",x"1e",x"d8",x"1e"),
  1301 => (x"e2",x"81",x"c8",x"49"),
  1302 => (x"86",x"c8",x"87",x"e2"),
  1303 => (x"48",x"66",x"c0",x"c1"),
  1304 => (x"c7",x"01",x"a8",x"c0"),
  1305 => (x"48",x"a6",x"c8",x"87"),
  1306 => (x"87",x"ce",x"78",x"c1"),
  1307 => (x"48",x"66",x"c0",x"c1"),
  1308 => (x"a6",x"d0",x"88",x"c1"),
  1309 => (x"e1",x"87",x"c3",x"58"),
  1310 => (x"a6",x"d0",x"87",x"ee"),
  1311 => (x"74",x"78",x"c2",x"48"),
  1312 => (x"cf",x"cd",x"02",x"9c"),
  1313 => (x"48",x"66",x"c8",x"87"),
  1314 => (x"a8",x"66",x"c4",x"c1"),
  1315 => (x"87",x"c4",x"cd",x"03"),
  1316 => (x"c0",x"48",x"a6",x"dc"),
  1317 => (x"c0",x"80",x"e8",x"78"),
  1318 => (x"87",x"dc",x"e0",x"78"),
  1319 => (x"d0",x"c1",x"4c",x"70"),
  1320 => (x"d7",x"c2",x"05",x"ac"),
  1321 => (x"7e",x"66",x"c4",x"87"),
  1322 => (x"c8",x"87",x"c0",x"e3"),
  1323 => (x"c7",x"e0",x"58",x"a6"),
  1324 => (x"c0",x"4c",x"70",x"87"),
  1325 => (x"c1",x"05",x"ac",x"ec"),
  1326 => (x"66",x"c8",x"87",x"ed"),
  1327 => (x"c0",x"91",x"cb",x"49"),
  1328 => (x"c4",x"81",x"66",x"fc"),
  1329 => (x"4d",x"6a",x"4a",x"a1"),
  1330 => (x"c4",x"4a",x"a1",x"c8"),
  1331 => (x"c3",x"c1",x"52",x"66"),
  1332 => (x"df",x"ff",x"79",x"dd"),
  1333 => (x"4c",x"70",x"87",x"e2"),
  1334 => (x"87",x"d9",x"02",x"9c"),
  1335 => (x"02",x"ac",x"fb",x"c0"),
  1336 => (x"55",x"74",x"87",x"d3"),
  1337 => (x"87",x"d0",x"df",x"ff"),
  1338 => (x"02",x"9c",x"4c",x"70"),
  1339 => (x"fb",x"c0",x"87",x"c7"),
  1340 => (x"ed",x"ff",x"05",x"ac"),
  1341 => (x"55",x"e0",x"c0",x"87"),
  1342 => (x"c0",x"55",x"c1",x"c2"),
  1343 => (x"66",x"d8",x"7d",x"97"),
  1344 => (x"05",x"a8",x"6e",x"48"),
  1345 => (x"66",x"c8",x"87",x"db"),
  1346 => (x"a8",x"66",x"cc",x"48"),
  1347 => (x"c8",x"87",x"ca",x"04"),
  1348 => (x"80",x"c1",x"48",x"66"),
  1349 => (x"c8",x"58",x"a6",x"cc"),
  1350 => (x"48",x"66",x"cc",x"87"),
  1351 => (x"a6",x"d0",x"88",x"c1"),
  1352 => (x"d3",x"de",x"ff",x"58"),
  1353 => (x"c1",x"4c",x"70",x"87"),
  1354 => (x"c8",x"05",x"ac",x"d0"),
  1355 => (x"48",x"66",x"d4",x"87"),
  1356 => (x"a6",x"d8",x"80",x"c1"),
  1357 => (x"ac",x"d0",x"c1",x"58"),
  1358 => (x"87",x"e9",x"fd",x"02"),
  1359 => (x"d8",x"48",x"66",x"c4"),
  1360 => (x"c9",x"05",x"a8",x"66"),
  1361 => (x"e0",x"c0",x"87",x"e0"),
  1362 => (x"78",x"c0",x"48",x"a6"),
  1363 => (x"fb",x"c0",x"48",x"74"),
  1364 => (x"48",x"7e",x"70",x"88"),
  1365 => (x"e2",x"c9",x"02",x"98"),
  1366 => (x"88",x"cb",x"48",x"87"),
  1367 => (x"98",x"48",x"7e",x"70"),
  1368 => (x"87",x"cd",x"c1",x"02"),
  1369 => (x"70",x"88",x"c9",x"48"),
  1370 => (x"02",x"98",x"48",x"7e"),
  1371 => (x"48",x"87",x"fe",x"c3"),
  1372 => (x"7e",x"70",x"88",x"c4"),
  1373 => (x"ce",x"02",x"98",x"48"),
  1374 => (x"88",x"c1",x"48",x"87"),
  1375 => (x"98",x"48",x"7e",x"70"),
  1376 => (x"87",x"e9",x"c3",x"02"),
  1377 => (x"dc",x"87",x"d6",x"c8"),
  1378 => (x"f0",x"c0",x"48",x"a6"),
  1379 => (x"e7",x"dc",x"ff",x"78"),
  1380 => (x"c0",x"4c",x"70",x"87"),
  1381 => (x"c0",x"02",x"ac",x"ec"),
  1382 => (x"e0",x"c0",x"87",x"c4"),
  1383 => (x"ec",x"c0",x"5c",x"a6"),
  1384 => (x"87",x"cd",x"02",x"ac"),
  1385 => (x"87",x"d0",x"dc",x"ff"),
  1386 => (x"ec",x"c0",x"4c",x"70"),
  1387 => (x"f3",x"ff",x"05",x"ac"),
  1388 => (x"ac",x"ec",x"c0",x"87"),
  1389 => (x"87",x"c4",x"c0",x"02"),
  1390 => (x"87",x"fc",x"db",x"ff"),
  1391 => (x"1e",x"ca",x"1e",x"c0"),
  1392 => (x"cb",x"49",x"66",x"d0"),
  1393 => (x"66",x"c4",x"c1",x"91"),
  1394 => (x"cc",x"80",x"71",x"48"),
  1395 => (x"66",x"c8",x"58",x"a6"),
  1396 => (x"d0",x"80",x"c4",x"48"),
  1397 => (x"66",x"cc",x"58",x"a6"),
  1398 => (x"dc",x"ff",x"49",x"bf"),
  1399 => (x"1e",x"c1",x"87",x"de"),
  1400 => (x"66",x"d4",x"1e",x"de"),
  1401 => (x"dc",x"ff",x"49",x"bf"),
  1402 => (x"86",x"d0",x"87",x"d2"),
  1403 => (x"c0",x"48",x"49",x"70"),
  1404 => (x"e8",x"c0",x"88",x"08"),
  1405 => (x"a8",x"c0",x"58",x"a6"),
  1406 => (x"87",x"ee",x"c0",x"06"),
  1407 => (x"48",x"66",x"e4",x"c0"),
  1408 => (x"c0",x"03",x"a8",x"dd"),
  1409 => (x"66",x"c4",x"87",x"e4"),
  1410 => (x"e4",x"c0",x"49",x"bf"),
  1411 => (x"e0",x"c0",x"81",x"66"),
  1412 => (x"66",x"e4",x"c0",x"51"),
  1413 => (x"c4",x"81",x"c1",x"49"),
  1414 => (x"c2",x"81",x"bf",x"66"),
  1415 => (x"e4",x"c0",x"51",x"c1"),
  1416 => (x"81",x"c2",x"49",x"66"),
  1417 => (x"81",x"bf",x"66",x"c4"),
  1418 => (x"48",x"6e",x"51",x"c0"),
  1419 => (x"78",x"ed",x"c9",x"c1"),
  1420 => (x"81",x"c8",x"49",x"6e"),
  1421 => (x"6e",x"51",x"66",x"d0"),
  1422 => (x"d4",x"81",x"c9",x"49"),
  1423 => (x"49",x"6e",x"51",x"66"),
  1424 => (x"66",x"dc",x"81",x"ca"),
  1425 => (x"48",x"66",x"d0",x"51"),
  1426 => (x"a6",x"d4",x"80",x"c1"),
  1427 => (x"48",x"66",x"c8",x"58"),
  1428 => (x"04",x"a8",x"66",x"cc"),
  1429 => (x"c8",x"87",x"cb",x"c0"),
  1430 => (x"80",x"c1",x"48",x"66"),
  1431 => (x"c5",x"58",x"a6",x"cc"),
  1432 => (x"66",x"cc",x"87",x"d9"),
  1433 => (x"d0",x"88",x"c1",x"48"),
  1434 => (x"ce",x"c5",x"58",x"a6"),
  1435 => (x"fa",x"db",x"ff",x"87"),
  1436 => (x"a6",x"e8",x"c0",x"87"),
  1437 => (x"f2",x"db",x"ff",x"58"),
  1438 => (x"a6",x"e0",x"c0",x"87"),
  1439 => (x"a8",x"ec",x"c0",x"58"),
  1440 => (x"87",x"ca",x"c0",x"05"),
  1441 => (x"c0",x"48",x"a6",x"dc"),
  1442 => (x"c0",x"78",x"66",x"e4"),
  1443 => (x"d8",x"ff",x"87",x"c4"),
  1444 => (x"66",x"c8",x"87",x"e6"),
  1445 => (x"c0",x"91",x"cb",x"49"),
  1446 => (x"71",x"48",x"66",x"fc"),
  1447 => (x"4a",x"7e",x"70",x"80"),
  1448 => (x"49",x"6e",x"82",x"c8"),
  1449 => (x"e4",x"c0",x"81",x"ca"),
  1450 => (x"66",x"dc",x"51",x"66"),
  1451 => (x"c0",x"81",x"c1",x"49"),
  1452 => (x"c1",x"89",x"66",x"e4"),
  1453 => (x"70",x"30",x"71",x"48"),
  1454 => (x"71",x"89",x"c1",x"49"),
  1455 => (x"ec",x"c2",x"7a",x"97"),
  1456 => (x"c0",x"49",x"bf",x"dc"),
  1457 => (x"97",x"29",x"66",x"e4"),
  1458 => (x"71",x"48",x"4a",x"6a"),
  1459 => (x"a6",x"ec",x"c0",x"98"),
  1460 => (x"c4",x"49",x"6e",x"58"),
  1461 => (x"d8",x"4d",x"69",x"81"),
  1462 => (x"66",x"c4",x"48",x"66"),
  1463 => (x"c8",x"c0",x"02",x"a8"),
  1464 => (x"48",x"a6",x"c4",x"87"),
  1465 => (x"c5",x"c0",x"78",x"c0"),
  1466 => (x"48",x"a6",x"c4",x"87"),
  1467 => (x"66",x"c4",x"78",x"c1"),
  1468 => (x"1e",x"e0",x"c0",x"1e"),
  1469 => (x"d8",x"ff",x"49",x"75"),
  1470 => (x"86",x"c8",x"87",x"c2"),
  1471 => (x"b7",x"c0",x"4c",x"70"),
  1472 => (x"d4",x"c1",x"06",x"ac"),
  1473 => (x"c0",x"85",x"74",x"87"),
  1474 => (x"89",x"74",x"49",x"e0"),
  1475 => (x"e0",x"c1",x"4b",x"75"),
  1476 => (x"fe",x"71",x"4a",x"d6"),
  1477 => (x"c2",x"87",x"d0",x"e6"),
  1478 => (x"66",x"e0",x"c0",x"85"),
  1479 => (x"c0",x"80",x"c1",x"48"),
  1480 => (x"c0",x"58",x"a6",x"e4"),
  1481 => (x"c1",x"49",x"66",x"e8"),
  1482 => (x"02",x"a9",x"70",x"81"),
  1483 => (x"c4",x"87",x"c8",x"c0"),
  1484 => (x"78",x"c0",x"48",x"a6"),
  1485 => (x"c4",x"87",x"c5",x"c0"),
  1486 => (x"78",x"c1",x"48",x"a6"),
  1487 => (x"c2",x"1e",x"66",x"c4"),
  1488 => (x"e0",x"c0",x"49",x"a4"),
  1489 => (x"70",x"88",x"71",x"48"),
  1490 => (x"49",x"75",x"1e",x"49"),
  1491 => (x"87",x"ec",x"d6",x"ff"),
  1492 => (x"b7",x"c0",x"86",x"c8"),
  1493 => (x"c0",x"ff",x"01",x"a8"),
  1494 => (x"66",x"e0",x"c0",x"87"),
  1495 => (x"87",x"d1",x"c0",x"02"),
  1496 => (x"81",x"c9",x"49",x"6e"),
  1497 => (x"51",x"66",x"e0",x"c0"),
  1498 => (x"ca",x"c1",x"48",x"6e"),
  1499 => (x"cc",x"c0",x"78",x"ee"),
  1500 => (x"c9",x"49",x"6e",x"87"),
  1501 => (x"6e",x"51",x"c2",x"81"),
  1502 => (x"da",x"cc",x"c1",x"48"),
  1503 => (x"48",x"66",x"c8",x"78"),
  1504 => (x"04",x"a8",x"66",x"cc"),
  1505 => (x"c8",x"87",x"cb",x"c0"),
  1506 => (x"80",x"c1",x"48",x"66"),
  1507 => (x"c0",x"58",x"a6",x"cc"),
  1508 => (x"66",x"cc",x"87",x"e9"),
  1509 => (x"d0",x"88",x"c1",x"48"),
  1510 => (x"de",x"c0",x"58",x"a6"),
  1511 => (x"c7",x"d5",x"ff",x"87"),
  1512 => (x"c0",x"4c",x"70",x"87"),
  1513 => (x"c6",x"c1",x"87",x"d5"),
  1514 => (x"c8",x"c0",x"05",x"ac"),
  1515 => (x"48",x"66",x"d0",x"87"),
  1516 => (x"a6",x"d4",x"80",x"c1"),
  1517 => (x"ef",x"d4",x"ff",x"58"),
  1518 => (x"d4",x"4c",x"70",x"87"),
  1519 => (x"80",x"c1",x"48",x"66"),
  1520 => (x"74",x"58",x"a6",x"d8"),
  1521 => (x"cb",x"c0",x"02",x"9c"),
  1522 => (x"48",x"66",x"c8",x"87"),
  1523 => (x"a8",x"66",x"c4",x"c1"),
  1524 => (x"87",x"fc",x"f2",x"04"),
  1525 => (x"87",x"c7",x"d4",x"ff"),
  1526 => (x"c7",x"48",x"66",x"c8"),
  1527 => (x"e5",x"c0",x"03",x"a8"),
  1528 => (x"f0",x"e8",x"c2",x"87"),
  1529 => (x"c8",x"78",x"c0",x"48"),
  1530 => (x"91",x"cb",x"49",x"66"),
  1531 => (x"81",x"66",x"fc",x"c0"),
  1532 => (x"6a",x"4a",x"a1",x"c4"),
  1533 => (x"79",x"52",x"c0",x"4a"),
  1534 => (x"c1",x"48",x"66",x"c8"),
  1535 => (x"58",x"a6",x"cc",x"80"),
  1536 => (x"ff",x"04",x"a8",x"c7"),
  1537 => (x"d4",x"ff",x"87",x"db"),
  1538 => (x"d6",x"de",x"ff",x"8e"),
  1539 => (x"61",x"6f",x"4c",x"87"),
  1540 => (x"2e",x"2a",x"20",x"64"),
  1541 => (x"20",x"3a",x"00",x"20"),
  1542 => (x"1e",x"73",x"1e",x"00"),
  1543 => (x"02",x"9b",x"4b",x"71"),
  1544 => (x"e8",x"c2",x"87",x"c6"),
  1545 => (x"78",x"c0",x"48",x"ec"),
  1546 => (x"e8",x"c2",x"1e",x"c7"),
  1547 => (x"c1",x"1e",x"bf",x"ec"),
  1548 => (x"c2",x"1e",x"e9",x"e4"),
  1549 => (x"49",x"bf",x"d4",x"e8"),
  1550 => (x"cc",x"87",x"ff",x"ed"),
  1551 => (x"d4",x"e8",x"c2",x"86"),
  1552 => (x"f7",x"e2",x"49",x"bf"),
  1553 => (x"02",x"9b",x"73",x"87"),
  1554 => (x"e4",x"c1",x"87",x"c8"),
  1555 => (x"e3",x"c0",x"49",x"e9"),
  1556 => (x"dd",x"ff",x"87",x"e2"),
  1557 => (x"73",x"1e",x"87",x"d1"),
  1558 => (x"c1",x"4b",x"c0",x"1e"),
  1559 => (x"c0",x"48",x"d5",x"e4"),
  1560 => (x"cc",x"e6",x"c1",x"50"),
  1561 => (x"d8",x"ff",x"49",x"bf"),
  1562 => (x"98",x"70",x"87",x"cd"),
  1563 => (x"c1",x"87",x"c4",x"05"),
  1564 => (x"73",x"4b",x"f9",x"e1"),
  1565 => (x"ee",x"dc",x"ff",x"48"),
  1566 => (x"4d",x"4f",x"52",x"87"),
  1567 => (x"61",x"6f",x"6c",x"20"),
  1568 => (x"67",x"6e",x"69",x"64"),
  1569 => (x"69",x"61",x"66",x"20"),
  1570 => (x"00",x"64",x"65",x"6c"),
  1571 => (x"87",x"e3",x"c7",x"1e"),
  1572 => (x"c4",x"fe",x"49",x"c1"),
  1573 => (x"fe",x"e8",x"fe",x"87"),
  1574 => (x"02",x"98",x"70",x"87"),
  1575 => (x"f1",x"fe",x"87",x"cd"),
  1576 => (x"98",x"70",x"87",x"f8"),
  1577 => (x"c1",x"87",x"c4",x"02"),
  1578 => (x"c0",x"87",x"c2",x"4a"),
  1579 => (x"05",x"9a",x"72",x"4a"),
  1580 => (x"1e",x"c0",x"87",x"ce"),
  1581 => (x"49",x"dc",x"e3",x"c1"),
  1582 => (x"87",x"ee",x"ee",x"c0"),
  1583 => (x"87",x"fe",x"86",x"c4"),
  1584 => (x"e3",x"c1",x"1e",x"c0"),
  1585 => (x"ee",x"c0",x"49",x"e7"),
  1586 => (x"1e",x"c0",x"87",x"e0"),
  1587 => (x"70",x"87",x"c7",x"fe"),
  1588 => (x"d5",x"ee",x"c0",x"49"),
  1589 => (x"87",x"da",x"c3",x"87"),
  1590 => (x"4f",x"26",x"8e",x"f8"),
  1591 => (x"66",x"20",x"44",x"53"),
  1592 => (x"65",x"6c",x"69",x"61"),
  1593 => (x"42",x"00",x"2e",x"64"),
  1594 => (x"69",x"74",x"6f",x"6f"),
  1595 => (x"2e",x"2e",x"67",x"6e"),
  1596 => (x"c0",x"1e",x"00",x"2e"),
  1597 => (x"c0",x"87",x"fa",x"e5"),
  1598 => (x"f6",x"87",x"e9",x"f1"),
  1599 => (x"1e",x"4f",x"26",x"87"),
  1600 => (x"48",x"ec",x"e8",x"c2"),
  1601 => (x"e8",x"c2",x"78",x"c0"),
  1602 => (x"78",x"c0",x"48",x"d4"),
  1603 => (x"e1",x"87",x"fd",x"fd"),
  1604 => (x"26",x"48",x"c0",x"87"),
  1605 => (x"01",x"00",x"00",x"4f"),
  1606 => (x"80",x"00",x"00",x"00"),
  1607 => (x"69",x"78",x"45",x"20"),
  1608 => (x"20",x"80",x"00",x"74"),
  1609 => (x"6b",x"63",x"61",x"42"),
  1610 => (x"00",x"10",x"2a",x"00"),
  1611 => (x"00",x"2a",x"40",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"00",x"10",x"2a"),
  1614 => (x"00",x"00",x"2a",x"5e"),
  1615 => (x"2a",x"00",x"00",x"00"),
  1616 => (x"7c",x"00",x"00",x"10"),
  1617 => (x"00",x"00",x"00",x"2a"),
  1618 => (x"10",x"2a",x"00",x"00"),
  1619 => (x"2a",x"9a",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"10",x"2a",x"00"),
  1622 => (x"00",x"2a",x"b8",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"00",x"10",x"2a"),
  1625 => (x"00",x"00",x"2a",x"d6"),
  1626 => (x"2a",x"00",x"00",x"00"),
  1627 => (x"f4",x"00",x"00",x"10"),
  1628 => (x"00",x"00",x"00",x"2a"),
  1629 => (x"10",x"dd",x"00",x"00"),
  1630 => (x"00",x"00",x"00",x"00"),
  1631 => (x"00",x"00",x"00",x"00"),
  1632 => (x"00",x"13",x"2b",x"00"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"00",x"00",x"19",x"90"),
  1636 => (x"39",x"39",x"49",x"54"),
  1637 => (x"20",x"20",x"41",x"34"),
  1638 => (x"00",x"4d",x"4f",x"52"),
  1639 => (x"48",x"f0",x"fe",x"1e"),
  1640 => (x"09",x"cd",x"78",x"c0"),
  1641 => (x"4f",x"26",x"09",x"79"),
  1642 => (x"f0",x"fe",x"1e",x"1e"),
  1643 => (x"26",x"48",x"7e",x"bf"),
  1644 => (x"fe",x"1e",x"4f",x"26"),
  1645 => (x"78",x"c1",x"48",x"f0"),
  1646 => (x"fe",x"1e",x"4f",x"26"),
  1647 => (x"78",x"c0",x"48",x"f0"),
  1648 => (x"71",x"1e",x"4f",x"26"),
  1649 => (x"52",x"52",x"c0",x"4a"),
  1650 => (x"5e",x"0e",x"4f",x"26"),
  1651 => (x"0e",x"5d",x"5c",x"5b"),
  1652 => (x"4d",x"71",x"86",x"f4"),
  1653 => (x"c1",x"7e",x"6d",x"97"),
  1654 => (x"6c",x"97",x"4c",x"a5"),
  1655 => (x"58",x"a6",x"c8",x"48"),
  1656 => (x"66",x"c4",x"48",x"6e"),
  1657 => (x"87",x"c5",x"05",x"a8"),
  1658 => (x"e6",x"c0",x"48",x"ff"),
  1659 => (x"87",x"ca",x"ff",x"87"),
  1660 => (x"97",x"49",x"a5",x"c2"),
  1661 => (x"a3",x"71",x"4b",x"6c"),
  1662 => (x"4b",x"6b",x"97",x"4b"),
  1663 => (x"6e",x"7e",x"6c",x"97"),
  1664 => (x"c8",x"80",x"c1",x"48"),
  1665 => (x"98",x"c7",x"58",x"a6"),
  1666 => (x"70",x"58",x"a6",x"cc"),
  1667 => (x"e1",x"fe",x"7c",x"97"),
  1668 => (x"f4",x"48",x"73",x"87"),
  1669 => (x"26",x"4d",x"26",x"8e"),
  1670 => (x"26",x"4b",x"26",x"4c"),
  1671 => (x"5b",x"5e",x"0e",x"4f"),
  1672 => (x"86",x"f4",x"0e",x"5c"),
  1673 => (x"66",x"d8",x"4c",x"71"),
  1674 => (x"9a",x"ff",x"c3",x"4a"),
  1675 => (x"97",x"4b",x"a4",x"c2"),
  1676 => (x"a1",x"73",x"49",x"6c"),
  1677 => (x"97",x"51",x"72",x"49"),
  1678 => (x"48",x"6e",x"7e",x"6c"),
  1679 => (x"a6",x"c8",x"80",x"c1"),
  1680 => (x"cc",x"98",x"c7",x"58"),
  1681 => (x"54",x"70",x"58",x"a6"),
  1682 => (x"ca",x"ff",x"8e",x"f4"),
  1683 => (x"fd",x"1e",x"1e",x"87"),
  1684 => (x"bf",x"e0",x"87",x"e8"),
  1685 => (x"e0",x"c0",x"49",x"4a"),
  1686 => (x"cb",x"02",x"99",x"c0"),
  1687 => (x"c2",x"1e",x"72",x"87"),
  1688 => (x"fe",x"49",x"d2",x"ec"),
  1689 => (x"86",x"c4",x"87",x"f7"),
  1690 => (x"70",x"87",x"fd",x"fc"),
  1691 => (x"87",x"c2",x"fd",x"7e"),
  1692 => (x"1e",x"4f",x"26",x"26"),
  1693 => (x"49",x"d2",x"ec",x"c2"),
  1694 => (x"c1",x"87",x"c7",x"fd"),
  1695 => (x"fc",x"49",x"cd",x"e9"),
  1696 => (x"f7",x"c3",x"87",x"da"),
  1697 => (x"0e",x"4f",x"26",x"87"),
  1698 => (x"5d",x"5c",x"5b",x"5e"),
  1699 => (x"c2",x"4d",x"71",x"0e"),
  1700 => (x"fc",x"49",x"d2",x"ec"),
  1701 => (x"4b",x"70",x"87",x"f4"),
  1702 => (x"04",x"ab",x"b7",x"c0"),
  1703 => (x"c3",x"87",x"c2",x"c3"),
  1704 => (x"c9",x"05",x"ab",x"f0"),
  1705 => (x"eb",x"ed",x"c1",x"87"),
  1706 => (x"c2",x"78",x"c1",x"48"),
  1707 => (x"e0",x"c3",x"87",x"e3"),
  1708 => (x"87",x"c9",x"05",x"ab"),
  1709 => (x"48",x"ef",x"ed",x"c1"),
  1710 => (x"d4",x"c2",x"78",x"c1"),
  1711 => (x"ef",x"ed",x"c1",x"87"),
  1712 => (x"87",x"c6",x"02",x"bf"),
  1713 => (x"4c",x"a3",x"c0",x"c2"),
  1714 => (x"4c",x"73",x"87",x"c2"),
  1715 => (x"bf",x"eb",x"ed",x"c1"),
  1716 => (x"87",x"e0",x"c0",x"02"),
  1717 => (x"b7",x"c4",x"49",x"74"),
  1718 => (x"ef",x"c1",x"91",x"29"),
  1719 => (x"4a",x"74",x"81",x"cb"),
  1720 => (x"92",x"c2",x"9a",x"cf"),
  1721 => (x"30",x"72",x"48",x"c1"),
  1722 => (x"ba",x"ff",x"4a",x"70"),
  1723 => (x"98",x"69",x"48",x"72"),
  1724 => (x"87",x"db",x"79",x"70"),
  1725 => (x"b7",x"c4",x"49",x"74"),
  1726 => (x"ef",x"c1",x"91",x"29"),
  1727 => (x"4a",x"74",x"81",x"cb"),
  1728 => (x"92",x"c2",x"9a",x"cf"),
  1729 => (x"30",x"72",x"48",x"c3"),
  1730 => (x"69",x"48",x"4a",x"70"),
  1731 => (x"75",x"79",x"70",x"b0"),
  1732 => (x"f0",x"c0",x"05",x"9d"),
  1733 => (x"48",x"d0",x"ff",x"87"),
  1734 => (x"ff",x"78",x"e1",x"c8"),
  1735 => (x"78",x"c5",x"48",x"d4"),
  1736 => (x"bf",x"ef",x"ed",x"c1"),
  1737 => (x"c3",x"87",x"c3",x"02"),
  1738 => (x"ed",x"c1",x"78",x"e0"),
  1739 => (x"c6",x"02",x"bf",x"eb"),
  1740 => (x"48",x"d4",x"ff",x"87"),
  1741 => (x"ff",x"78",x"f0",x"c3"),
  1742 => (x"0b",x"7b",x"0b",x"d4"),
  1743 => (x"c8",x"48",x"d0",x"ff"),
  1744 => (x"e0",x"c0",x"78",x"e1"),
  1745 => (x"ef",x"ed",x"c1",x"78"),
  1746 => (x"c1",x"78",x"c0",x"48"),
  1747 => (x"c0",x"48",x"eb",x"ed"),
  1748 => (x"d2",x"ec",x"c2",x"78"),
  1749 => (x"87",x"f2",x"f9",x"49"),
  1750 => (x"b7",x"c0",x"4b",x"70"),
  1751 => (x"fe",x"fc",x"03",x"ab"),
  1752 => (x"26",x"48",x"c0",x"87"),
  1753 => (x"26",x"4c",x"26",x"4d"),
  1754 => (x"00",x"4f",x"26",x"4b"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"1e",x"00",x"00",x"00"),
  1757 => (x"fc",x"49",x"4a",x"71"),
  1758 => (x"4f",x"26",x"87",x"cd"),
  1759 => (x"72",x"4a",x"c0",x"1e"),
  1760 => (x"c1",x"91",x"c4",x"49"),
  1761 => (x"c0",x"81",x"cb",x"ef"),
  1762 => (x"d0",x"82",x"c1",x"79"),
  1763 => (x"ee",x"04",x"aa",x"b7"),
  1764 => (x"0e",x"4f",x"26",x"87"),
  1765 => (x"5d",x"5c",x"5b",x"5e"),
  1766 => (x"f8",x"4d",x"71",x"0e"),
  1767 => (x"4a",x"75",x"87",x"dc"),
  1768 => (x"92",x"2a",x"b7",x"c4"),
  1769 => (x"82",x"cb",x"ef",x"c1"),
  1770 => (x"9c",x"cf",x"4c",x"75"),
  1771 => (x"49",x"6a",x"94",x"c2"),
  1772 => (x"c3",x"2b",x"74",x"4b"),
  1773 => (x"74",x"48",x"c2",x"9b"),
  1774 => (x"ff",x"4c",x"70",x"30"),
  1775 => (x"71",x"48",x"74",x"bc"),
  1776 => (x"f7",x"7a",x"70",x"98"),
  1777 => (x"48",x"73",x"87",x"ec"),
  1778 => (x"00",x"87",x"d8",x"fe"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"1e",x"00",x"00",x"00"),
  1795 => (x"c8",x"48",x"d0",x"ff"),
  1796 => (x"48",x"71",x"78",x"e1"),
  1797 => (x"78",x"08",x"d4",x"ff"),
  1798 => (x"ff",x"1e",x"4f",x"26"),
  1799 => (x"e1",x"c8",x"48",x"d0"),
  1800 => (x"ff",x"48",x"71",x"78"),
  1801 => (x"c4",x"78",x"08",x"d4"),
  1802 => (x"d4",x"ff",x"48",x"66"),
  1803 => (x"4f",x"26",x"78",x"08"),
  1804 => (x"c4",x"4a",x"71",x"1e"),
  1805 => (x"72",x"1e",x"49",x"66"),
  1806 => (x"87",x"de",x"ff",x"49"),
  1807 => (x"c0",x"48",x"d0",x"ff"),
  1808 => (x"26",x"26",x"78",x"e0"),
  1809 => (x"1e",x"73",x"1e",x"4f"),
  1810 => (x"66",x"c8",x"4b",x"71"),
  1811 => (x"4a",x"73",x"1e",x"49"),
  1812 => (x"49",x"a2",x"e0",x"c1"),
  1813 => (x"26",x"87",x"d9",x"ff"),
  1814 => (x"4d",x"26",x"87",x"c4"),
  1815 => (x"4b",x"26",x"4c",x"26"),
  1816 => (x"ff",x"1e",x"4f",x"26"),
  1817 => (x"ff",x"c3",x"4a",x"d4"),
  1818 => (x"48",x"d0",x"ff",x"7a"),
  1819 => (x"de",x"78",x"e1",x"c0"),
  1820 => (x"dc",x"ec",x"c2",x"7a"),
  1821 => (x"48",x"49",x"7a",x"bf"),
  1822 => (x"7a",x"70",x"28",x"c8"),
  1823 => (x"28",x"d0",x"48",x"71"),
  1824 => (x"48",x"71",x"7a",x"70"),
  1825 => (x"7a",x"70",x"28",x"d8"),
  1826 => (x"c0",x"48",x"d0",x"ff"),
  1827 => (x"4f",x"26",x"78",x"e0"),
  1828 => (x"48",x"d0",x"ff",x"1e"),
  1829 => (x"71",x"78",x"c9",x"c8"),
  1830 => (x"08",x"d4",x"ff",x"48"),
  1831 => (x"1e",x"4f",x"26",x"78"),
  1832 => (x"eb",x"49",x"4a",x"71"),
  1833 => (x"48",x"d0",x"ff",x"87"),
  1834 => (x"4f",x"26",x"78",x"c8"),
  1835 => (x"71",x"1e",x"73",x"1e"),
  1836 => (x"ec",x"ec",x"c2",x"4b"),
  1837 => (x"87",x"c3",x"02",x"bf"),
  1838 => (x"ff",x"87",x"eb",x"c2"),
  1839 => (x"c9",x"c8",x"48",x"d0"),
  1840 => (x"c0",x"48",x"73",x"78"),
  1841 => (x"d4",x"ff",x"b0",x"e0"),
  1842 => (x"ec",x"c2",x"78",x"08"),
  1843 => (x"78",x"c0",x"48",x"e0"),
  1844 => (x"c5",x"02",x"66",x"c8"),
  1845 => (x"49",x"ff",x"c3",x"87"),
  1846 => (x"49",x"c0",x"87",x"c2"),
  1847 => (x"59",x"e8",x"ec",x"c2"),
  1848 => (x"c6",x"02",x"66",x"cc"),
  1849 => (x"d5",x"d5",x"c5",x"87"),
  1850 => (x"cf",x"87",x"c4",x"4a"),
  1851 => (x"c2",x"4a",x"ff",x"ff"),
  1852 => (x"c2",x"5a",x"ec",x"ec"),
  1853 => (x"c1",x"48",x"ec",x"ec"),
  1854 => (x"26",x"87",x"c4",x"78"),
  1855 => (x"26",x"4c",x"26",x"4d"),
  1856 => (x"0e",x"4f",x"26",x"4b"),
  1857 => (x"5d",x"5c",x"5b",x"5e"),
  1858 => (x"c2",x"4a",x"71",x"0e"),
  1859 => (x"4c",x"bf",x"e8",x"ec"),
  1860 => (x"cb",x"02",x"9a",x"72"),
  1861 => (x"91",x"c8",x"49",x"87"),
  1862 => (x"4b",x"e2",x"f2",x"c1"),
  1863 => (x"87",x"c4",x"83",x"71"),
  1864 => (x"4b",x"e2",x"f6",x"c1"),
  1865 => (x"49",x"13",x"4d",x"c0"),
  1866 => (x"ec",x"c2",x"99",x"74"),
  1867 => (x"71",x"48",x"bf",x"e4"),
  1868 => (x"08",x"d4",x"ff",x"b8"),
  1869 => (x"2c",x"b7",x"c1",x"78"),
  1870 => (x"ad",x"b7",x"c8",x"85"),
  1871 => (x"c2",x"87",x"e7",x"04"),
  1872 => (x"48",x"bf",x"e0",x"ec"),
  1873 => (x"ec",x"c2",x"80",x"c8"),
  1874 => (x"ee",x"fe",x"58",x"e4"),
  1875 => (x"1e",x"73",x"1e",x"87"),
  1876 => (x"4a",x"13",x"4b",x"71"),
  1877 => (x"87",x"cb",x"02",x"9a"),
  1878 => (x"e6",x"fe",x"49",x"72"),
  1879 => (x"9a",x"4a",x"13",x"87"),
  1880 => (x"fe",x"87",x"f5",x"05"),
  1881 => (x"c2",x"1e",x"87",x"d9"),
  1882 => (x"49",x"bf",x"e0",x"ec"),
  1883 => (x"48",x"e0",x"ec",x"c2"),
  1884 => (x"c4",x"78",x"a1",x"c1"),
  1885 => (x"03",x"a9",x"b7",x"c0"),
  1886 => (x"d4",x"ff",x"87",x"db"),
  1887 => (x"e4",x"ec",x"c2",x"48"),
  1888 => (x"ec",x"c2",x"78",x"bf"),
  1889 => (x"c2",x"49",x"bf",x"e0"),
  1890 => (x"c1",x"48",x"e0",x"ec"),
  1891 => (x"c0",x"c4",x"78",x"a1"),
  1892 => (x"e5",x"04",x"a9",x"b7"),
  1893 => (x"48",x"d0",x"ff",x"87"),
  1894 => (x"ec",x"c2",x"78",x"c8"),
  1895 => (x"78",x"c0",x"48",x"ec"),
  1896 => (x"00",x"00",x"4f",x"26"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"5f",x"5f",x"00"),
  1900 => (x"03",x"00",x"00",x"00"),
  1901 => (x"03",x"03",x"00",x"03"),
  1902 => (x"7f",x"14",x"00",x"00"),
  1903 => (x"7f",x"7f",x"14",x"7f"),
  1904 => (x"24",x"00",x"00",x"14"),
  1905 => (x"3a",x"6b",x"6b",x"2e"),
  1906 => (x"6a",x"4c",x"00",x"12"),
  1907 => (x"56",x"6c",x"18",x"36"),
  1908 => (x"7e",x"30",x"00",x"32"),
  1909 => (x"3a",x"77",x"59",x"4f"),
  1910 => (x"00",x"00",x"40",x"68"),
  1911 => (x"00",x"03",x"07",x"04"),
  1912 => (x"00",x"00",x"00",x"00"),
  1913 => (x"41",x"63",x"3e",x"1c"),
  1914 => (x"00",x"00",x"00",x"00"),
  1915 => (x"1c",x"3e",x"63",x"41"),
  1916 => (x"2a",x"08",x"00",x"00"),
  1917 => (x"3e",x"1c",x"1c",x"3e"),
  1918 => (x"08",x"00",x"08",x"2a"),
  1919 => (x"08",x"3e",x"3e",x"08"),
  1920 => (x"00",x"00",x"00",x"08"),
  1921 => (x"00",x"60",x"e0",x"80"),
  1922 => (x"08",x"00",x"00",x"00"),
  1923 => (x"08",x"08",x"08",x"08"),
  1924 => (x"00",x"00",x"00",x"08"),
  1925 => (x"00",x"60",x"60",x"00"),
  1926 => (x"60",x"40",x"00",x"00"),
  1927 => (x"06",x"0c",x"18",x"30"),
  1928 => (x"3e",x"00",x"01",x"03"),
  1929 => (x"7f",x"4d",x"59",x"7f"),
  1930 => (x"04",x"00",x"00",x"3e"),
  1931 => (x"00",x"7f",x"7f",x"06"),
  1932 => (x"42",x"00",x"00",x"00"),
  1933 => (x"4f",x"59",x"71",x"63"),
  1934 => (x"22",x"00",x"00",x"46"),
  1935 => (x"7f",x"49",x"49",x"63"),
  1936 => (x"1c",x"18",x"00",x"36"),
  1937 => (x"7f",x"7f",x"13",x"16"),
  1938 => (x"27",x"00",x"00",x"10"),
  1939 => (x"7d",x"45",x"45",x"67"),
  1940 => (x"3c",x"00",x"00",x"39"),
  1941 => (x"79",x"49",x"4b",x"7e"),
  1942 => (x"01",x"00",x"00",x"30"),
  1943 => (x"0f",x"79",x"71",x"01"),
  1944 => (x"36",x"00",x"00",x"07"),
  1945 => (x"7f",x"49",x"49",x"7f"),
  1946 => (x"06",x"00",x"00",x"36"),
  1947 => (x"3f",x"69",x"49",x"4f"),
  1948 => (x"00",x"00",x"00",x"1e"),
  1949 => (x"00",x"66",x"66",x"00"),
  1950 => (x"00",x"00",x"00",x"00"),
  1951 => (x"00",x"66",x"e6",x"80"),
  1952 => (x"08",x"00",x"00",x"00"),
  1953 => (x"22",x"14",x"14",x"08"),
  1954 => (x"14",x"00",x"00",x"22"),
  1955 => (x"14",x"14",x"14",x"14"),
  1956 => (x"22",x"00",x"00",x"14"),
  1957 => (x"08",x"14",x"14",x"22"),
  1958 => (x"02",x"00",x"00",x"08"),
  1959 => (x"0f",x"59",x"51",x"03"),
  1960 => (x"7f",x"3e",x"00",x"06"),
  1961 => (x"1f",x"55",x"5d",x"41"),
  1962 => (x"7e",x"00",x"00",x"1e"),
  1963 => (x"7f",x"09",x"09",x"7f"),
  1964 => (x"7f",x"00",x"00",x"7e"),
  1965 => (x"7f",x"49",x"49",x"7f"),
  1966 => (x"1c",x"00",x"00",x"36"),
  1967 => (x"41",x"41",x"63",x"3e"),
  1968 => (x"7f",x"00",x"00",x"41"),
  1969 => (x"3e",x"63",x"41",x"7f"),
  1970 => (x"7f",x"00",x"00",x"1c"),
  1971 => (x"41",x"49",x"49",x"7f"),
  1972 => (x"7f",x"00",x"00",x"41"),
  1973 => (x"01",x"09",x"09",x"7f"),
  1974 => (x"3e",x"00",x"00",x"01"),
  1975 => (x"7b",x"49",x"41",x"7f"),
  1976 => (x"7f",x"00",x"00",x"7a"),
  1977 => (x"7f",x"08",x"08",x"7f"),
  1978 => (x"00",x"00",x"00",x"7f"),
  1979 => (x"41",x"7f",x"7f",x"41"),
  1980 => (x"20",x"00",x"00",x"00"),
  1981 => (x"7f",x"40",x"40",x"60"),
  1982 => (x"7f",x"7f",x"00",x"3f"),
  1983 => (x"63",x"36",x"1c",x"08"),
  1984 => (x"7f",x"00",x"00",x"41"),
  1985 => (x"40",x"40",x"40",x"7f"),
  1986 => (x"7f",x"7f",x"00",x"40"),
  1987 => (x"7f",x"06",x"0c",x"06"),
  1988 => (x"7f",x"7f",x"00",x"7f"),
  1989 => (x"7f",x"18",x"0c",x"06"),
  1990 => (x"3e",x"00",x"00",x"7f"),
  1991 => (x"7f",x"41",x"41",x"7f"),
  1992 => (x"7f",x"00",x"00",x"3e"),
  1993 => (x"0f",x"09",x"09",x"7f"),
  1994 => (x"7f",x"3e",x"00",x"06"),
  1995 => (x"7e",x"7f",x"61",x"41"),
  1996 => (x"7f",x"00",x"00",x"40"),
  1997 => (x"7f",x"19",x"09",x"7f"),
  1998 => (x"26",x"00",x"00",x"66"),
  1999 => (x"7b",x"59",x"4d",x"6f"),
  2000 => (x"01",x"00",x"00",x"32"),
  2001 => (x"01",x"7f",x"7f",x"01"),
  2002 => (x"3f",x"00",x"00",x"01"),
  2003 => (x"7f",x"40",x"40",x"7f"),
  2004 => (x"0f",x"00",x"00",x"3f"),
  2005 => (x"3f",x"70",x"70",x"3f"),
  2006 => (x"7f",x"7f",x"00",x"0f"),
  2007 => (x"7f",x"30",x"18",x"30"),
  2008 => (x"63",x"41",x"00",x"7f"),
  2009 => (x"36",x"1c",x"1c",x"36"),
  2010 => (x"03",x"01",x"41",x"63"),
  2011 => (x"06",x"7c",x"7c",x"06"),
  2012 => (x"71",x"61",x"01",x"03"),
  2013 => (x"43",x"47",x"4d",x"59"),
  2014 => (x"00",x"00",x"00",x"41"),
  2015 => (x"41",x"41",x"7f",x"7f"),
  2016 => (x"03",x"01",x"00",x"00"),
  2017 => (x"30",x"18",x"0c",x"06"),
  2018 => (x"00",x"00",x"40",x"60"),
  2019 => (x"7f",x"7f",x"41",x"41"),
  2020 => (x"0c",x"08",x"00",x"00"),
  2021 => (x"0c",x"06",x"03",x"06"),
  2022 => (x"80",x"80",x"00",x"08"),
  2023 => (x"80",x"80",x"80",x"80"),
  2024 => (x"00",x"00",x"00",x"80"),
  2025 => (x"04",x"07",x"03",x"00"),
  2026 => (x"20",x"00",x"00",x"00"),
  2027 => (x"7c",x"54",x"54",x"74"),
  2028 => (x"7f",x"00",x"00",x"78"),
  2029 => (x"7c",x"44",x"44",x"7f"),
  2030 => (x"38",x"00",x"00",x"38"),
  2031 => (x"44",x"44",x"44",x"7c"),
  2032 => (x"38",x"00",x"00",x"00"),
  2033 => (x"7f",x"44",x"44",x"7c"),
  2034 => (x"38",x"00",x"00",x"7f"),
  2035 => (x"5c",x"54",x"54",x"7c"),
  2036 => (x"04",x"00",x"00",x"18"),
  2037 => (x"05",x"05",x"7f",x"7e"),
  2038 => (x"18",x"00",x"00",x"00"),
  2039 => (x"fc",x"a4",x"a4",x"bc"),
  2040 => (x"7f",x"00",x"00",x"7c"),
  2041 => (x"7c",x"04",x"04",x"7f"),
  2042 => (x"00",x"00",x"00",x"78"),
  2043 => (x"40",x"7d",x"3d",x"00"),
  2044 => (x"80",x"00",x"00",x"00"),
  2045 => (x"7d",x"fd",x"80",x"80"),
  2046 => (x"7f",x"00",x"00",x"00"),
  2047 => (x"6c",x"38",x"10",x"7f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

