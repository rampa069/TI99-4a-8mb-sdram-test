
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"00",x"44"),
     1 => (x"40",x"7f",x"3f",x"00"),
     2 => (x"7c",x"7c",x"00",x"00"),
     3 => (x"7c",x"0c",x"18",x"0c"),
     4 => (x"7c",x"00",x"00",x"78"),
     5 => (x"7c",x"04",x"04",x"7c"),
     6 => (x"38",x"00",x"00",x"78"),
     7 => (x"7c",x"44",x"44",x"7c"),
     8 => (x"fc",x"00",x"00",x"38"),
     9 => (x"3c",x"24",x"24",x"fc"),
    10 => (x"18",x"00",x"00",x"18"),
    11 => (x"fc",x"24",x"24",x"3c"),
    12 => (x"7c",x"00",x"00",x"fc"),
    13 => (x"0c",x"04",x"04",x"7c"),
    14 => (x"48",x"00",x"00",x"08"),
    15 => (x"74",x"54",x"54",x"5c"),
    16 => (x"04",x"00",x"00",x"20"),
    17 => (x"44",x"44",x"7f",x"3f"),
    18 => (x"3c",x"00",x"00",x"00"),
    19 => (x"7c",x"40",x"40",x"7c"),
    20 => (x"1c",x"00",x"00",x"7c"),
    21 => (x"3c",x"60",x"60",x"3c"),
    22 => (x"7c",x"3c",x"00",x"1c"),
    23 => (x"7c",x"60",x"30",x"60"),
    24 => (x"6c",x"44",x"00",x"3c"),
    25 => (x"6c",x"38",x"10",x"38"),
    26 => (x"1c",x"00",x"00",x"44"),
    27 => (x"3c",x"60",x"e0",x"bc"),
    28 => (x"44",x"00",x"00",x"1c"),
    29 => (x"4c",x"5c",x"74",x"64"),
    30 => (x"08",x"00",x"00",x"44"),
    31 => (x"41",x"77",x"3e",x"08"),
    32 => (x"00",x"00",x"00",x"41"),
    33 => (x"00",x"7f",x"7f",x"00"),
    34 => (x"41",x"00",x"00",x"00"),
    35 => (x"08",x"3e",x"77",x"41"),
    36 => (x"01",x"02",x"00",x"08"),
    37 => (x"02",x"02",x"03",x"01"),
    38 => (x"7f",x"7f",x"00",x"01"),
    39 => (x"7f",x"7f",x"7f",x"7f"),
    40 => (x"08",x"08",x"00",x"7f"),
    41 => (x"3e",x"3e",x"1c",x"1c"),
    42 => (x"7f",x"7f",x"7f",x"7f"),
    43 => (x"1c",x"1c",x"3e",x"3e"),
    44 => (x"10",x"00",x"08",x"08"),
    45 => (x"18",x"7c",x"7c",x"18"),
    46 => (x"10",x"00",x"00",x"10"),
    47 => (x"30",x"7c",x"7c",x"30"),
    48 => (x"30",x"10",x"00",x"10"),
    49 => (x"1e",x"78",x"60",x"60"),
    50 => (x"66",x"42",x"00",x"06"),
    51 => (x"66",x"3c",x"18",x"3c"),
    52 => (x"38",x"78",x"00",x"42"),
    53 => (x"6c",x"c6",x"c2",x"6a"),
    54 => (x"00",x"60",x"00",x"38"),
    55 => (x"00",x"00",x"60",x"00"),
    56 => (x"5e",x"0e",x"00",x"60"),
    57 => (x"0e",x"5d",x"5c",x"5b"),
    58 => (x"c2",x"4c",x"71",x"1e"),
    59 => (x"4d",x"bf",x"fd",x"ec"),
    60 => (x"1e",x"c0",x"4b",x"c0"),
    61 => (x"c7",x"02",x"ab",x"74"),
    62 => (x"48",x"a6",x"c4",x"87"),
    63 => (x"87",x"c5",x"78",x"c0"),
    64 => (x"c1",x"48",x"a6",x"c4"),
    65 => (x"1e",x"66",x"c4",x"78"),
    66 => (x"df",x"ee",x"49",x"73"),
    67 => (x"c0",x"86",x"c8",x"87"),
    68 => (x"ee",x"ef",x"49",x"e0"),
    69 => (x"4a",x"a5",x"c4",x"87"),
    70 => (x"f0",x"f0",x"49",x"6a"),
    71 => (x"87",x"c6",x"f1",x"87"),
    72 => (x"83",x"c1",x"85",x"cb"),
    73 => (x"04",x"ab",x"b7",x"c8"),
    74 => (x"26",x"87",x"c7",x"ff"),
    75 => (x"4c",x"26",x"4d",x"26"),
    76 => (x"4f",x"26",x"4b",x"26"),
    77 => (x"c2",x"4a",x"71",x"1e"),
    78 => (x"c2",x"5a",x"c1",x"ed"),
    79 => (x"c7",x"48",x"c1",x"ed"),
    80 => (x"dd",x"fe",x"49",x"78"),
    81 => (x"1e",x"4f",x"26",x"87"),
    82 => (x"4a",x"71",x"1e",x"73"),
    83 => (x"03",x"aa",x"b7",x"c0"),
    84 => (x"d3",x"c2",x"87",x"d3"),
    85 => (x"c4",x"05",x"bf",x"c3"),
    86 => (x"c2",x"4b",x"c1",x"87"),
    87 => (x"c2",x"4b",x"c0",x"87"),
    88 => (x"c4",x"5b",x"c7",x"d3"),
    89 => (x"c7",x"d3",x"c2",x"87"),
    90 => (x"c3",x"d3",x"c2",x"5a"),
    91 => (x"9a",x"c1",x"4a",x"bf"),
    92 => (x"49",x"a2",x"c0",x"c1"),
    93 => (x"fc",x"87",x"e8",x"ec"),
    94 => (x"c3",x"d3",x"c2",x"48"),
    95 => (x"ef",x"fe",x"78",x"bf"),
    96 => (x"4a",x"71",x"1e",x"87"),
    97 => (x"72",x"1e",x"66",x"c4"),
    98 => (x"87",x"f9",x"ea",x"49"),
    99 => (x"1e",x"4f",x"26",x"26"),
   100 => (x"c3",x"48",x"d4",x"ff"),
   101 => (x"d0",x"ff",x"78",x"ff"),
   102 => (x"78",x"e1",x"c0",x"48"),
   103 => (x"c1",x"48",x"d4",x"ff"),
   104 => (x"c4",x"48",x"71",x"78"),
   105 => (x"08",x"d4",x"ff",x"30"),
   106 => (x"48",x"d0",x"ff",x"78"),
   107 => (x"26",x"78",x"e0",x"c0"),
   108 => (x"d3",x"c2",x"1e",x"4f"),
   109 => (x"e6",x"49",x"bf",x"c3"),
   110 => (x"ec",x"c2",x"87",x"f9"),
   111 => (x"bf",x"e8",x"48",x"f5"),
   112 => (x"f1",x"ec",x"c2",x"78"),
   113 => (x"78",x"bf",x"ec",x"48"),
   114 => (x"bf",x"f5",x"ec",x"c2"),
   115 => (x"ff",x"c3",x"49",x"4a"),
   116 => (x"2a",x"b7",x"c8",x"99"),
   117 => (x"b0",x"71",x"48",x"72"),
   118 => (x"58",x"fd",x"ec",x"c2"),
   119 => (x"5e",x"0e",x"4f",x"26"),
   120 => (x"0e",x"5d",x"5c",x"5b"),
   121 => (x"c8",x"ff",x"4b",x"71"),
   122 => (x"f0",x"ec",x"c2",x"87"),
   123 => (x"73",x"50",x"c0",x"48"),
   124 => (x"87",x"df",x"e6",x"49"),
   125 => (x"c2",x"4c",x"49",x"70"),
   126 => (x"49",x"ee",x"cb",x"9c"),
   127 => (x"70",x"87",x"cc",x"cb"),
   128 => (x"f0",x"ec",x"c2",x"4d"),
   129 => (x"c1",x"05",x"bf",x"97"),
   130 => (x"66",x"d0",x"87",x"e2"),
   131 => (x"f9",x"ec",x"c2",x"49"),
   132 => (x"d6",x"05",x"99",x"bf"),
   133 => (x"49",x"66",x"d4",x"87"),
   134 => (x"bf",x"f1",x"ec",x"c2"),
   135 => (x"87",x"cb",x"05",x"99"),
   136 => (x"ee",x"e5",x"49",x"73"),
   137 => (x"02",x"98",x"70",x"87"),
   138 => (x"c1",x"87",x"c1",x"c1"),
   139 => (x"87",x"c1",x"fe",x"4c"),
   140 => (x"e2",x"ca",x"49",x"75"),
   141 => (x"02",x"98",x"70",x"87"),
   142 => (x"ec",x"c2",x"87",x"c6"),
   143 => (x"50",x"c1",x"48",x"f0"),
   144 => (x"97",x"f0",x"ec",x"c2"),
   145 => (x"e3",x"c0",x"05",x"bf"),
   146 => (x"f9",x"ec",x"c2",x"87"),
   147 => (x"66",x"d0",x"49",x"bf"),
   148 => (x"d6",x"ff",x"05",x"99"),
   149 => (x"f1",x"ec",x"c2",x"87"),
   150 => (x"66",x"d4",x"49",x"bf"),
   151 => (x"ca",x"ff",x"05",x"99"),
   152 => (x"e4",x"49",x"73",x"87"),
   153 => (x"98",x"70",x"87",x"ed"),
   154 => (x"87",x"ff",x"fe",x"05"),
   155 => (x"fb",x"fa",x"48",x"74"),
   156 => (x"5b",x"5e",x"0e",x"87"),
   157 => (x"f8",x"0e",x"5d",x"5c"),
   158 => (x"4c",x"4d",x"c0",x"86"),
   159 => (x"c4",x"7e",x"bf",x"ec"),
   160 => (x"ec",x"c2",x"48",x"a6"),
   161 => (x"c1",x"78",x"bf",x"fd"),
   162 => (x"c7",x"1e",x"c0",x"1e"),
   163 => (x"87",x"ce",x"fd",x"49"),
   164 => (x"98",x"70",x"86",x"c8"),
   165 => (x"ff",x"87",x"cd",x"02"),
   166 => (x"87",x"eb",x"fa",x"49"),
   167 => (x"e3",x"49",x"da",x"c1"),
   168 => (x"4d",x"c1",x"87",x"f1"),
   169 => (x"97",x"f0",x"ec",x"c2"),
   170 => (x"87",x"cf",x"02",x"bf"),
   171 => (x"bf",x"fb",x"d2",x"c2"),
   172 => (x"c2",x"b9",x"c1",x"49"),
   173 => (x"71",x"59",x"ff",x"d2"),
   174 => (x"c2",x"87",x"d4",x"fb"),
   175 => (x"4b",x"bf",x"f5",x"ec"),
   176 => (x"bf",x"c3",x"d3",x"c2"),
   177 => (x"87",x"e9",x"c0",x"05"),
   178 => (x"e3",x"49",x"fd",x"c3"),
   179 => (x"fa",x"c3",x"87",x"c5"),
   180 => (x"87",x"ff",x"e2",x"49"),
   181 => (x"ff",x"c3",x"49",x"73"),
   182 => (x"c0",x"1e",x"71",x"99"),
   183 => (x"87",x"e1",x"fa",x"49"),
   184 => (x"b7",x"c8",x"49",x"73"),
   185 => (x"c1",x"1e",x"71",x"29"),
   186 => (x"87",x"d5",x"fa",x"49"),
   187 => (x"f4",x"c5",x"86",x"c8"),
   188 => (x"f9",x"ec",x"c2",x"87"),
   189 => (x"02",x"9b",x"4b",x"bf"),
   190 => (x"d2",x"c2",x"87",x"dd"),
   191 => (x"c7",x"49",x"bf",x"ff"),
   192 => (x"98",x"70",x"87",x"d5"),
   193 => (x"c0",x"87",x"c4",x"05"),
   194 => (x"c2",x"87",x"d2",x"4b"),
   195 => (x"fa",x"c6",x"49",x"e0"),
   196 => (x"c3",x"d3",x"c2",x"87"),
   197 => (x"c2",x"87",x"c6",x"58"),
   198 => (x"c0",x"48",x"ff",x"d2"),
   199 => (x"c2",x"49",x"73",x"78"),
   200 => (x"87",x"cd",x"05",x"99"),
   201 => (x"e1",x"49",x"eb",x"c3"),
   202 => (x"49",x"70",x"87",x"e9"),
   203 => (x"c2",x"02",x"99",x"c2"),
   204 => (x"73",x"4c",x"fb",x"87"),
   205 => (x"05",x"99",x"c1",x"49"),
   206 => (x"f4",x"c3",x"87",x"cd"),
   207 => (x"87",x"d3",x"e1",x"49"),
   208 => (x"99",x"c2",x"49",x"70"),
   209 => (x"fa",x"87",x"c2",x"02"),
   210 => (x"c8",x"49",x"73",x"4c"),
   211 => (x"87",x"cd",x"05",x"99"),
   212 => (x"e0",x"49",x"f5",x"c3"),
   213 => (x"49",x"70",x"87",x"fd"),
   214 => (x"d5",x"02",x"99",x"c2"),
   215 => (x"c1",x"ed",x"c2",x"87"),
   216 => (x"87",x"ca",x"02",x"bf"),
   217 => (x"c2",x"88",x"c1",x"48"),
   218 => (x"c0",x"58",x"c5",x"ed"),
   219 => (x"4c",x"ff",x"87",x"c2"),
   220 => (x"49",x"73",x"4d",x"c1"),
   221 => (x"cd",x"05",x"99",x"c4"),
   222 => (x"49",x"f2",x"c3",x"87"),
   223 => (x"70",x"87",x"d4",x"e0"),
   224 => (x"02",x"99",x"c2",x"49"),
   225 => (x"ed",x"c2",x"87",x"dc"),
   226 => (x"48",x"7e",x"bf",x"c1"),
   227 => (x"03",x"a8",x"b7",x"c7"),
   228 => (x"6e",x"87",x"cb",x"c0"),
   229 => (x"c2",x"80",x"c1",x"48"),
   230 => (x"c0",x"58",x"c5",x"ed"),
   231 => (x"4c",x"fe",x"87",x"c2"),
   232 => (x"fd",x"c3",x"4d",x"c1"),
   233 => (x"ea",x"df",x"ff",x"49"),
   234 => (x"c2",x"49",x"70",x"87"),
   235 => (x"87",x"d5",x"02",x"99"),
   236 => (x"bf",x"c1",x"ed",x"c2"),
   237 => (x"87",x"c9",x"c0",x"02"),
   238 => (x"48",x"c1",x"ed",x"c2"),
   239 => (x"c2",x"c0",x"78",x"c0"),
   240 => (x"c1",x"4c",x"fd",x"87"),
   241 => (x"49",x"fa",x"c3",x"4d"),
   242 => (x"87",x"c7",x"df",x"ff"),
   243 => (x"99",x"c2",x"49",x"70"),
   244 => (x"87",x"d9",x"c0",x"02"),
   245 => (x"bf",x"c1",x"ed",x"c2"),
   246 => (x"a8",x"b7",x"c7",x"48"),
   247 => (x"87",x"c9",x"c0",x"03"),
   248 => (x"48",x"c1",x"ed",x"c2"),
   249 => (x"c2",x"c0",x"78",x"c7"),
   250 => (x"c1",x"4c",x"fc",x"87"),
   251 => (x"ac",x"b7",x"c0",x"4d"),
   252 => (x"87",x"d3",x"c0",x"03"),
   253 => (x"c1",x"48",x"66",x"c4"),
   254 => (x"7e",x"70",x"80",x"d8"),
   255 => (x"c0",x"02",x"bf",x"6e"),
   256 => (x"74",x"4b",x"87",x"c5"),
   257 => (x"c0",x"0f",x"73",x"49"),
   258 => (x"1e",x"f0",x"c3",x"1e"),
   259 => (x"f7",x"49",x"da",x"c1"),
   260 => (x"86",x"c8",x"87",x"cc"),
   261 => (x"c0",x"02",x"98",x"70"),
   262 => (x"ed",x"c2",x"87",x"d8"),
   263 => (x"6e",x"7e",x"bf",x"c1"),
   264 => (x"c4",x"91",x"cb",x"49"),
   265 => (x"82",x"71",x"4a",x"66"),
   266 => (x"c5",x"c0",x"02",x"6a"),
   267 => (x"49",x"6e",x"4b",x"87"),
   268 => (x"9d",x"75",x"0f",x"73"),
   269 => (x"87",x"c8",x"c0",x"02"),
   270 => (x"bf",x"c1",x"ed",x"c2"),
   271 => (x"87",x"e2",x"f2",x"49"),
   272 => (x"bf",x"c7",x"d3",x"c2"),
   273 => (x"87",x"dd",x"c0",x"02"),
   274 => (x"87",x"cb",x"c2",x"49"),
   275 => (x"c0",x"02",x"98",x"70"),
   276 => (x"ed",x"c2",x"87",x"d3"),
   277 => (x"f2",x"49",x"bf",x"c1"),
   278 => (x"49",x"c0",x"87",x"c8"),
   279 => (x"c2",x"87",x"e8",x"f3"),
   280 => (x"c0",x"48",x"c7",x"d3"),
   281 => (x"f3",x"8e",x"f8",x"78"),
   282 => (x"5e",x"0e",x"87",x"c2"),
   283 => (x"0e",x"5d",x"5c",x"5b"),
   284 => (x"c2",x"4c",x"71",x"1e"),
   285 => (x"49",x"bf",x"fd",x"ec"),
   286 => (x"4d",x"a1",x"cd",x"c1"),
   287 => (x"69",x"81",x"d1",x"c1"),
   288 => (x"02",x"9c",x"74",x"7e"),
   289 => (x"a5",x"c4",x"87",x"cf"),
   290 => (x"c2",x"7b",x"74",x"4b"),
   291 => (x"49",x"bf",x"fd",x"ec"),
   292 => (x"6e",x"87",x"e1",x"f2"),
   293 => (x"05",x"9c",x"74",x"7b"),
   294 => (x"4b",x"c0",x"87",x"c4"),
   295 => (x"4b",x"c1",x"87",x"c2"),
   296 => (x"e2",x"f2",x"49",x"73"),
   297 => (x"02",x"66",x"d4",x"87"),
   298 => (x"de",x"49",x"87",x"c7"),
   299 => (x"c2",x"4a",x"70",x"87"),
   300 => (x"c2",x"4a",x"c0",x"87"),
   301 => (x"26",x"5a",x"cb",x"d3"),
   302 => (x"00",x"87",x"f1",x"f1"),
   303 => (x"00",x"00",x"00",x"00"),
   304 => (x"00",x"00",x"00",x"00"),
   305 => (x"00",x"00",x"00",x"00"),
   306 => (x"1e",x"00",x"00",x"00"),
   307 => (x"c8",x"ff",x"4a",x"71"),
   308 => (x"a1",x"72",x"49",x"bf"),
   309 => (x"1e",x"4f",x"26",x"48"),
   310 => (x"89",x"bf",x"c8",x"ff"),
   311 => (x"c0",x"c0",x"c0",x"fe"),
   312 => (x"01",x"a9",x"c0",x"c0"),
   313 => (x"4a",x"c0",x"87",x"c4"),
   314 => (x"4a",x"c1",x"87",x"c2"),
   315 => (x"4f",x"26",x"48",x"72"),
   316 => (x"5c",x"5b",x"5e",x"0e"),
   317 => (x"4b",x"71",x"0e",x"5d"),
   318 => (x"d0",x"4c",x"d4",x"ff"),
   319 => (x"78",x"c0",x"48",x"66"),
   320 => (x"dc",x"ff",x"49",x"d6"),
   321 => (x"ff",x"c3",x"87",x"c5"),
   322 => (x"c3",x"49",x"6c",x"7c"),
   323 => (x"4d",x"71",x"99",x"ff"),
   324 => (x"99",x"f0",x"c3",x"49"),
   325 => (x"05",x"a9",x"e0",x"c1"),
   326 => (x"ff",x"c3",x"87",x"cb"),
   327 => (x"c3",x"48",x"6c",x"7c"),
   328 => (x"08",x"66",x"d0",x"98"),
   329 => (x"7c",x"ff",x"c3",x"78"),
   330 => (x"c8",x"49",x"4a",x"6c"),
   331 => (x"7c",x"ff",x"c3",x"31"),
   332 => (x"b2",x"71",x"4a",x"6c"),
   333 => (x"31",x"c8",x"49",x"72"),
   334 => (x"6c",x"7c",x"ff",x"c3"),
   335 => (x"72",x"b2",x"71",x"4a"),
   336 => (x"c3",x"31",x"c8",x"49"),
   337 => (x"4a",x"6c",x"7c",x"ff"),
   338 => (x"d0",x"ff",x"b2",x"71"),
   339 => (x"78",x"e0",x"c0",x"48"),
   340 => (x"c2",x"02",x"9b",x"73"),
   341 => (x"75",x"7b",x"72",x"87"),
   342 => (x"26",x"4d",x"26",x"48"),
   343 => (x"26",x"4b",x"26",x"4c"),
   344 => (x"4f",x"26",x"1e",x"4f"),
   345 => (x"5c",x"5b",x"5e",x"0e"),
   346 => (x"76",x"86",x"f8",x"0e"),
   347 => (x"49",x"a6",x"c8",x"1e"),
   348 => (x"c4",x"87",x"fd",x"fd"),
   349 => (x"6e",x"4b",x"70",x"86"),
   350 => (x"03",x"a8",x"c4",x"48"),
   351 => (x"73",x"87",x"f0",x"c2"),
   352 => (x"9a",x"f0",x"c3",x"4a"),
   353 => (x"02",x"aa",x"d0",x"c1"),
   354 => (x"e0",x"c1",x"87",x"c7"),
   355 => (x"de",x"c2",x"05",x"aa"),
   356 => (x"c8",x"49",x"73",x"87"),
   357 => (x"87",x"c3",x"02",x"99"),
   358 => (x"73",x"87",x"c6",x"ff"),
   359 => (x"c2",x"9c",x"c3",x"4c"),
   360 => (x"c2",x"c1",x"05",x"ac"),
   361 => (x"49",x"66",x"c4",x"87"),
   362 => (x"1e",x"71",x"31",x"c9"),
   363 => (x"d4",x"4a",x"66",x"c4"),
   364 => (x"c5",x"ed",x"c2",x"92"),
   365 => (x"fe",x"81",x"72",x"49"),
   366 => (x"d8",x"87",x"ce",x"d0"),
   367 => (x"ca",x"d9",x"ff",x"49"),
   368 => (x"1e",x"c0",x"c8",x"87"),
   369 => (x"49",x"e2",x"db",x"c2"),
   370 => (x"87",x"d2",x"ec",x"fd"),
   371 => (x"c0",x"48",x"d0",x"ff"),
   372 => (x"db",x"c2",x"78",x"e0"),
   373 => (x"66",x"cc",x"1e",x"e2"),
   374 => (x"c2",x"92",x"d4",x"4a"),
   375 => (x"72",x"49",x"c5",x"ed"),
   376 => (x"d6",x"ce",x"fe",x"81"),
   377 => (x"c1",x"86",x"cc",x"87"),
   378 => (x"c2",x"c1",x"05",x"ac"),
   379 => (x"49",x"66",x"c4",x"87"),
   380 => (x"1e",x"71",x"31",x"c9"),
   381 => (x"d4",x"4a",x"66",x"c4"),
   382 => (x"c5",x"ed",x"c2",x"92"),
   383 => (x"fe",x"81",x"72",x"49"),
   384 => (x"c2",x"87",x"c6",x"cf"),
   385 => (x"c8",x"1e",x"e2",x"db"),
   386 => (x"92",x"d4",x"4a",x"66"),
   387 => (x"49",x"c5",x"ed",x"c2"),
   388 => (x"cc",x"fe",x"81",x"72"),
   389 => (x"49",x"d7",x"87",x"d7"),
   390 => (x"87",x"ef",x"d7",x"ff"),
   391 => (x"c2",x"1e",x"c0",x"c8"),
   392 => (x"fd",x"49",x"e2",x"db"),
   393 => (x"cc",x"87",x"d0",x"ea"),
   394 => (x"48",x"d0",x"ff",x"86"),
   395 => (x"f8",x"78",x"e0",x"c0"),
   396 => (x"87",x"e7",x"fc",x"8e"),
   397 => (x"5c",x"5b",x"5e",x"0e"),
   398 => (x"71",x"1e",x"0e",x"5d"),
   399 => (x"4c",x"d4",x"ff",x"4d"),
   400 => (x"48",x"7e",x"66",x"d4"),
   401 => (x"06",x"a8",x"b7",x"c3"),
   402 => (x"48",x"c0",x"87",x"c5"),
   403 => (x"75",x"87",x"e9",x"c1"),
   404 => (x"fe",x"dc",x"fe",x"49"),
   405 => (x"c4",x"1e",x"75",x"87"),
   406 => (x"93",x"d4",x"4b",x"66"),
   407 => (x"83",x"c5",x"ed",x"c2"),
   408 => (x"c6",x"fe",x"49",x"73"),
   409 => (x"83",x"c8",x"87",x"d3"),
   410 => (x"d0",x"ff",x"4b",x"6b"),
   411 => (x"78",x"e1",x"c8",x"48"),
   412 => (x"48",x"73",x"7c",x"dd"),
   413 => (x"70",x"98",x"ff",x"c3"),
   414 => (x"c8",x"49",x"73",x"7c"),
   415 => (x"48",x"71",x"29",x"b7"),
   416 => (x"70",x"98",x"ff",x"c3"),
   417 => (x"d0",x"49",x"73",x"7c"),
   418 => (x"48",x"71",x"29",x"b7"),
   419 => (x"70",x"98",x"ff",x"c3"),
   420 => (x"d8",x"48",x"73",x"7c"),
   421 => (x"7c",x"70",x"28",x"b7"),
   422 => (x"7c",x"7c",x"7c",x"c0"),
   423 => (x"7c",x"7c",x"7c",x"7c"),
   424 => (x"7c",x"7c",x"7c",x"7c"),
   425 => (x"48",x"d0",x"ff",x"7c"),
   426 => (x"c4",x"78",x"e0",x"c0"),
   427 => (x"49",x"dc",x"1e",x"66"),
   428 => (x"87",x"fc",x"d5",x"ff"),
   429 => (x"48",x"73",x"86",x"c8"),
   430 => (x"87",x"dd",x"fa",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

