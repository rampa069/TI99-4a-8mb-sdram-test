library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00000044",
     1 => x"407f3f00",
     2 => x"7c7c0000",
     3 => x"7c0c180c",
     4 => x"7c000078",
     5 => x"7c04047c",
     6 => x"38000078",
     7 => x"7c44447c",
     8 => x"fc000038",
     9 => x"3c2424fc",
    10 => x"18000018",
    11 => x"fc24243c",
    12 => x"7c0000fc",
    13 => x"0c04047c",
    14 => x"48000008",
    15 => x"7454545c",
    16 => x"04000020",
    17 => x"44447f3f",
    18 => x"3c000000",
    19 => x"7c40407c",
    20 => x"1c00007c",
    21 => x"3c60603c",
    22 => x"7c3c001c",
    23 => x"7c603060",
    24 => x"6c44003c",
    25 => x"6c381038",
    26 => x"1c000044",
    27 => x"3c60e0bc",
    28 => x"4400001c",
    29 => x"4c5c7464",
    30 => x"08000044",
    31 => x"41773e08",
    32 => x"00000041",
    33 => x"007f7f00",
    34 => x"41000000",
    35 => x"083e7741",
    36 => x"01020008",
    37 => x"02020301",
    38 => x"7f7f0001",
    39 => x"7f7f7f7f",
    40 => x"0808007f",
    41 => x"3e3e1c1c",
    42 => x"7f7f7f7f",
    43 => x"1c1c3e3e",
    44 => x"10000808",
    45 => x"187c7c18",
    46 => x"10000010",
    47 => x"307c7c30",
    48 => x"30100010",
    49 => x"1e786060",
    50 => x"66420006",
    51 => x"663c183c",
    52 => x"38780042",
    53 => x"6cc6c26a",
    54 => x"00600038",
    55 => x"00006000",
    56 => x"5e0e0060",
    57 => x"0e5d5c5b",
    58 => x"c24c711e",
    59 => x"4dbffdec",
    60 => x"1ec04bc0",
    61 => x"c702ab74",
    62 => x"48a6c487",
    63 => x"87c578c0",
    64 => x"c148a6c4",
    65 => x"1e66c478",
    66 => x"dfee4973",
    67 => x"c086c887",
    68 => x"eeef49e0",
    69 => x"4aa5c487",
    70 => x"f0f0496a",
    71 => x"87c6f187",
    72 => x"83c185cb",
    73 => x"04abb7c8",
    74 => x"2687c7ff",
    75 => x"4c264d26",
    76 => x"4f264b26",
    77 => x"c24a711e",
    78 => x"c25ac1ed",
    79 => x"c748c1ed",
    80 => x"ddfe4978",
    81 => x"1e4f2687",
    82 => x"4a711e73",
    83 => x"03aab7c0",
    84 => x"d3c287d3",
    85 => x"c405bfc3",
    86 => x"c24bc187",
    87 => x"c24bc087",
    88 => x"c45bc7d3",
    89 => x"c7d3c287",
    90 => x"c3d3c25a",
    91 => x"9ac14abf",
    92 => x"49a2c0c1",
    93 => x"fc87e8ec",
    94 => x"c3d3c248",
    95 => x"effe78bf",
    96 => x"4a711e87",
    97 => x"721e66c4",
    98 => x"87f9ea49",
    99 => x"1e4f2626",
   100 => x"c348d4ff",
   101 => x"d0ff78ff",
   102 => x"78e1c048",
   103 => x"c148d4ff",
   104 => x"c4487178",
   105 => x"08d4ff30",
   106 => x"48d0ff78",
   107 => x"2678e0c0",
   108 => x"d3c21e4f",
   109 => x"e649bfc3",
   110 => x"ecc287f9",
   111 => x"bfe848f5",
   112 => x"f1ecc278",
   113 => x"78bfec48",
   114 => x"bff5ecc2",
   115 => x"ffc3494a",
   116 => x"2ab7c899",
   117 => x"b0714872",
   118 => x"58fdecc2",
   119 => x"5e0e4f26",
   120 => x"0e5d5c5b",
   121 => x"c8ff4b71",
   122 => x"f0ecc287",
   123 => x"7350c048",
   124 => x"87dfe649",
   125 => x"c24c4970",
   126 => x"49eecb9c",
   127 => x"7087cccb",
   128 => x"f0ecc24d",
   129 => x"c105bf97",
   130 => x"66d087e2",
   131 => x"f9ecc249",
   132 => x"d60599bf",
   133 => x"4966d487",
   134 => x"bff1ecc2",
   135 => x"87cb0599",
   136 => x"eee54973",
   137 => x"02987087",
   138 => x"c187c1c1",
   139 => x"87c1fe4c",
   140 => x"e2ca4975",
   141 => x"02987087",
   142 => x"ecc287c6",
   143 => x"50c148f0",
   144 => x"97f0ecc2",
   145 => x"e3c005bf",
   146 => x"f9ecc287",
   147 => x"66d049bf",
   148 => x"d6ff0599",
   149 => x"f1ecc287",
   150 => x"66d449bf",
   151 => x"caff0599",
   152 => x"e4497387",
   153 => x"987087ed",
   154 => x"87fffe05",
   155 => x"fbfa4874",
   156 => x"5b5e0e87",
   157 => x"f80e5d5c",
   158 => x"4c4dc086",
   159 => x"c47ebfec",
   160 => x"ecc248a6",
   161 => x"c178bffd",
   162 => x"c71ec01e",
   163 => x"87cefd49",
   164 => x"987086c8",
   165 => x"ff87cd02",
   166 => x"87ebfa49",
   167 => x"e349dac1",
   168 => x"4dc187f1",
   169 => x"97f0ecc2",
   170 => x"87cf02bf",
   171 => x"bffbd2c2",
   172 => x"c2b9c149",
   173 => x"7159ffd2",
   174 => x"c287d4fb",
   175 => x"4bbff5ec",
   176 => x"bfc3d3c2",
   177 => x"87e9c005",
   178 => x"e349fdc3",
   179 => x"fac387c5",
   180 => x"87ffe249",
   181 => x"ffc34973",
   182 => x"c01e7199",
   183 => x"87e1fa49",
   184 => x"b7c84973",
   185 => x"c11e7129",
   186 => x"87d5fa49",
   187 => x"f4c586c8",
   188 => x"f9ecc287",
   189 => x"029b4bbf",
   190 => x"d2c287dd",
   191 => x"c749bfff",
   192 => x"987087d5",
   193 => x"c087c405",
   194 => x"c287d24b",
   195 => x"fac649e0",
   196 => x"c3d3c287",
   197 => x"c287c658",
   198 => x"c048ffd2",
   199 => x"c2497378",
   200 => x"87cd0599",
   201 => x"e149ebc3",
   202 => x"497087e9",
   203 => x"c20299c2",
   204 => x"734cfb87",
   205 => x"0599c149",
   206 => x"f4c387cd",
   207 => x"87d3e149",
   208 => x"99c24970",
   209 => x"fa87c202",
   210 => x"c849734c",
   211 => x"87cd0599",
   212 => x"e049f5c3",
   213 => x"497087fd",
   214 => x"d50299c2",
   215 => x"c1edc287",
   216 => x"87ca02bf",
   217 => x"c288c148",
   218 => x"c058c5ed",
   219 => x"4cff87c2",
   220 => x"49734dc1",
   221 => x"cd0599c4",
   222 => x"49f2c387",
   223 => x"7087d4e0",
   224 => x"0299c249",
   225 => x"edc287dc",
   226 => x"487ebfc1",
   227 => x"03a8b7c7",
   228 => x"6e87cbc0",
   229 => x"c280c148",
   230 => x"c058c5ed",
   231 => x"4cfe87c2",
   232 => x"fdc34dc1",
   233 => x"eadfff49",
   234 => x"c2497087",
   235 => x"87d50299",
   236 => x"bfc1edc2",
   237 => x"87c9c002",
   238 => x"48c1edc2",
   239 => x"c2c078c0",
   240 => x"c14cfd87",
   241 => x"49fac34d",
   242 => x"87c7dfff",
   243 => x"99c24970",
   244 => x"87d9c002",
   245 => x"bfc1edc2",
   246 => x"a8b7c748",
   247 => x"87c9c003",
   248 => x"48c1edc2",
   249 => x"c2c078c7",
   250 => x"c14cfc87",
   251 => x"acb7c04d",
   252 => x"87d3c003",
   253 => x"c14866c4",
   254 => x"7e7080d8",
   255 => x"c002bf6e",
   256 => x"744b87c5",
   257 => x"c00f7349",
   258 => x"1ef0c31e",
   259 => x"f749dac1",
   260 => x"86c887cc",
   261 => x"c0029870",
   262 => x"edc287d8",
   263 => x"6e7ebfc1",
   264 => x"c491cb49",
   265 => x"82714a66",
   266 => x"c5c0026a",
   267 => x"496e4b87",
   268 => x"9d750f73",
   269 => x"87c8c002",
   270 => x"bfc1edc2",
   271 => x"87e2f249",
   272 => x"bfc7d3c2",
   273 => x"87ddc002",
   274 => x"87cbc249",
   275 => x"c0029870",
   276 => x"edc287d3",
   277 => x"f249bfc1",
   278 => x"49c087c8",
   279 => x"c287e8f3",
   280 => x"c048c7d3",
   281 => x"f38ef878",
   282 => x"5e0e87c2",
   283 => x"0e5d5c5b",
   284 => x"c24c711e",
   285 => x"49bffdec",
   286 => x"4da1cdc1",
   287 => x"6981d1c1",
   288 => x"029c747e",
   289 => x"a5c487cf",
   290 => x"c27b744b",
   291 => x"49bffdec",
   292 => x"6e87e1f2",
   293 => x"059c747b",
   294 => x"4bc087c4",
   295 => x"4bc187c2",
   296 => x"e2f24973",
   297 => x"0266d487",
   298 => x"de4987c7",
   299 => x"c24a7087",
   300 => x"c24ac087",
   301 => x"265acbd3",
   302 => x"0087f1f1",
   303 => x"00000000",
   304 => x"00000000",
   305 => x"00000000",
   306 => x"1e000000",
   307 => x"c8ff4a71",
   308 => x"a17249bf",
   309 => x"1e4f2648",
   310 => x"89bfc8ff",
   311 => x"c0c0c0fe",
   312 => x"01a9c0c0",
   313 => x"4ac087c4",
   314 => x"4ac187c2",
   315 => x"4f264872",
   316 => x"5c5b5e0e",
   317 => x"4b710e5d",
   318 => x"d04cd4ff",
   319 => x"78c04866",
   320 => x"dcff49d6",
   321 => x"ffc387c5",
   322 => x"c3496c7c",
   323 => x"4d7199ff",
   324 => x"99f0c349",
   325 => x"05a9e0c1",
   326 => x"ffc387cb",
   327 => x"c3486c7c",
   328 => x"0866d098",
   329 => x"7cffc378",
   330 => x"c8494a6c",
   331 => x"7cffc331",
   332 => x"b2714a6c",
   333 => x"31c84972",
   334 => x"6c7cffc3",
   335 => x"72b2714a",
   336 => x"c331c849",
   337 => x"4a6c7cff",
   338 => x"d0ffb271",
   339 => x"78e0c048",
   340 => x"c2029b73",
   341 => x"757b7287",
   342 => x"264d2648",
   343 => x"264b264c",
   344 => x"4f261e4f",
   345 => x"5c5b5e0e",
   346 => x"7686f80e",
   347 => x"49a6c81e",
   348 => x"c487fdfd",
   349 => x"6e4b7086",
   350 => x"03a8c448",
   351 => x"7387f0c2",
   352 => x"9af0c34a",
   353 => x"02aad0c1",
   354 => x"e0c187c7",
   355 => x"dec205aa",
   356 => x"c8497387",
   357 => x"87c30299",
   358 => x"7387c6ff",
   359 => x"c29cc34c",
   360 => x"c2c105ac",
   361 => x"4966c487",
   362 => x"1e7131c9",
   363 => x"d44a66c4",
   364 => x"c5edc292",
   365 => x"fe817249",
   366 => x"d887ced0",
   367 => x"cad9ff49",
   368 => x"1ec0c887",
   369 => x"49e2dbc2",
   370 => x"87d2ecfd",
   371 => x"c048d0ff",
   372 => x"dbc278e0",
   373 => x"66cc1ee2",
   374 => x"c292d44a",
   375 => x"7249c5ed",
   376 => x"d6cefe81",
   377 => x"c186cc87",
   378 => x"c2c105ac",
   379 => x"4966c487",
   380 => x"1e7131c9",
   381 => x"d44a66c4",
   382 => x"c5edc292",
   383 => x"fe817249",
   384 => x"c287c6cf",
   385 => x"c81ee2db",
   386 => x"92d44a66",
   387 => x"49c5edc2",
   388 => x"ccfe8172",
   389 => x"49d787d7",
   390 => x"87efd7ff",
   391 => x"c21ec0c8",
   392 => x"fd49e2db",
   393 => x"cc87d0ea",
   394 => x"48d0ff86",
   395 => x"f878e0c0",
   396 => x"87e7fc8e",
   397 => x"5c5b5e0e",
   398 => x"711e0e5d",
   399 => x"4cd4ff4d",
   400 => x"487e66d4",
   401 => x"06a8b7c3",
   402 => x"48c087c5",
   403 => x"7587e9c1",
   404 => x"fedcfe49",
   405 => x"c41e7587",
   406 => x"93d44b66",
   407 => x"83c5edc2",
   408 => x"c6fe4973",
   409 => x"83c887d3",
   410 => x"d0ff4b6b",
   411 => x"78e1c848",
   412 => x"48737cdd",
   413 => x"7098ffc3",
   414 => x"c849737c",
   415 => x"487129b7",
   416 => x"7098ffc3",
   417 => x"d049737c",
   418 => x"487129b7",
   419 => x"7098ffc3",
   420 => x"d848737c",
   421 => x"7c7028b7",
   422 => x"7c7c7cc0",
   423 => x"7c7c7c7c",
   424 => x"7c7c7c7c",
   425 => x"48d0ff7c",
   426 => x"c478e0c0",
   427 => x"49dc1e66",
   428 => x"87fcd5ff",
   429 => x"487386c8",
   430 => x"87ddfa26",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
